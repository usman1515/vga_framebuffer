----------------------------------------------------------------------------------
-- Company:
-- Engineer:
--
-- Design Name:
-- Module Name: ram_init_phillips_pm5544_grayscale - Behavioral
-- Project Name:
-- Target Devices:
-- Tool Versions: 2021.2
-- Description:
--
-- Dependencies:
--
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
----------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;


package ram_init_phillips_pm5544_grayscale is

    constant FB_WIDTH : integer := 640;
    constant FB_HEIGHT : integer := 480;
    constant FB_PIXELS : integer := FB_WIDTH * FB_HEIGHT;

    constant DATA_WIDTH : integer := 4;
    constant DEPTH : integer := FB_PIXELS;

    subtype addr_t is integer range 0 to DEPTH - 1;
    subtype ram_word_t is std_logic_vector(DATA_WIDTH-1 downto 0);

    type ram_type is array (addr_t) of ram_word_t;

    -- Synthesizable constant RAM content
    constant INIT_RAM : ram_type := (
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"A",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"4",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"4",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"A",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"A",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"4",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"A",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"A",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"4",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"A",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"A",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"4",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"4",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"A",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"A",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"4",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"A",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"A",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"4",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"A",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"A",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"4",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"4",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"A",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"A",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"4",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"A",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"A",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"4",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"A",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"A",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"4",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"4",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"A",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"A",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"4",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"A",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"A",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"4",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"A",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"A",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"4",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"4",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"A",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"A",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"4",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"A",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"A",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"4",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"A",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"A",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",
        x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",
        x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",
        x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",
        x"2",    x"2",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"6",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",
        x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",
        x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",
        x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",
        x"2",    x"6",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",
        x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",
        x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",
        x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",
        x"2",    x"A",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"A",
        x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",
        x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",
        x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",
        x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",
        x"2",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"6",
        x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",
        x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",
        x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",
        x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",
        x"6",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"2",
        x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",
        x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",
        x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",
        x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",
        x"A",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"A",    x"2",
        x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",
        x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",
        x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",
        x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"6",    x"2",
        x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",
        x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",
        x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",
        x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"6",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"2",    x"2",
        x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",
        x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",
        x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",
        x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"A",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"D",    x"F",
        x"D",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"F",    x"F",    x"C",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"F",    x"F",
        x"B",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"B",    x"F",    x"F",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"C",    x"F",    x"F",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"D",    x"F",    x"E",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"E",    x"F",    x"D",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"F",    x"F",    x"C",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"F",    x"F",    x"B",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"B",    x"F",    x"F",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"C",    x"F",    x"F",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"D",    x"F",    x"E",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"E",    x"F",    x"D",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"F",    x"F",    x"C",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"F",    x"F",    x"B",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"B",
        x"F",    x"F",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"C",    x"F",    x"F",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"D",
        x"F",    x"D",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"8",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"8",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"8",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"8",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"8",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"8",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"8",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"8",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"8",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"8",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"8",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"8",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"8",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"8",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",
        x"8",    x"9",    x"A",    x"B",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"E",
        x"E",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"B",    x"A",    x"9",    x"8",
        x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"8",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"A",
        x"C",    x"D",    x"D",    x"E",    x"E",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"E",    x"E",    x"D",    x"D",    x"C",
        x"A",    x"9",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"8",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"A",
        x"C",    x"D",    x"D",    x"E",    x"E",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"E",    x"E",    x"D",    x"D",    x"C",
        x"A",    x"8",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"8",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"9",    x"B",    x"D",    x"E",    x"E",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"E",    x"E",    x"D",    x"C",    x"A",    x"8",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"8",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"B",    x"C",    x"E",    x"E",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"E",    x"E",    x"C",    x"B",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"8",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"9",
        x"C",    x"D",    x"E",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"E",    x"E",    x"C",
        x"A",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"8",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"F",    x"F",    x"C",    x"C",    x"E",    x"E",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"E",    x"D",    x"D",    x"F",    x"F",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"8",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"C",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"C",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"8",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"B",    x"D",    x"E",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"E",    x"E",    x"C",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"8",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"9",    x"C",    x"E",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"E",    x"D",    x"A",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"8",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"A",    x"D",    x"E",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"E",    x"D",    x"A",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"8",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"9",    x"D",    x"E",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"E",    x"D",    x"A",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"8",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"9",
        x"D",    x"E",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"E",    x"D",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"8",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"9",    x"D",    x"E",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"E",    x"D",    x"9",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"8",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"B",    x"E",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"E",    x"C",    x"8",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"8",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"9",
        x"D",    x"E",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"E",    x"D",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"8",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"8",    x"B",    x"E",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"E",    x"C",    x"8",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"8",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",
        x"7",    x"7",    x"9",    x"D",    x"E",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"E",    x"D",    x"9",    x"7",    x"7",
        x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"8",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"D",    x"F",
        x"D",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"F",    x"F",    x"C",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"F",    x"F",
        x"B",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"B",    x"F",    x"F",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"C",    x"F",    x"F",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"D",    x"F",    x"E",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"E",    x"F",    x"D",
        x"B",    x"E",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"E",    x"C",
        x"D",    x"F",    x"E",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"E",    x"F",    x"D",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"F",    x"F",    x"C",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"F",    x"F",    x"B",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"B",
        x"F",    x"F",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"C",    x"F",    x"F",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"D",
        x"F",    x"D",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"6",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"B",    x"F",    x"F",    x"9",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"B",    x"F",    x"F",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"C",    x"F",    x"E",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"9",    x"D",    x"E",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"6",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"E",    x"D",    x"9",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"E",    x"F",    x"C",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"F",    x"F",    x"B",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"9",    x"F",    x"F",    x"B",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"8",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"A",    x"F",    x"F",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"8",
        x"C",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"6",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"D",
        x"8",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"7",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"C",    x"E",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"6",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"D",    x"8",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"7",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"C",    x"E",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"6",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"E",    x"D",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"7",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"C",    x"E",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"6",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"E",    x"C",    x"8",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"7",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"E",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"6",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"E",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"7",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",    x"E",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"6",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"E",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"7",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"9",    x"E",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"6",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"E",    x"9",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"7",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"8",    x"D",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"6",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"D",    x"8",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"7",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"E",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"6",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"E",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"7",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"E",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"6",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"E",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"7",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"D",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"6",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"D",    x"8",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"7",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"B",    x"E",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"6",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"E",    x"B",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"7",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"8",    x"D",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"6",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"E",    x"8",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"7",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"B",    x"E",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"6",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"E",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"7",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"9",
        x"E",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"6",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"E",
        x"9",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"7",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"D",    x"7",    x"7",    x"C",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"6",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"C",    x"7",    x"7",    x"D",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"7",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"D",    x"8",    x"E",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"6",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"E",    x"8",    x"D",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"7",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"E",    x"E",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"6",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"E",    x"E",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"7",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"6",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"7",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"9",    x"E",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"6",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"E",    x"A",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"7",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"6",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"7",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"E",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"6",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"E",    x"8",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"7",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"A",    x"E",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"6",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"E",    x"A",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"7",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"C",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"6",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"C",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"7",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"D",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"6",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"D",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"7",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"9",    x"E",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"6",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"E",    x"9",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"7",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"E",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"6",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"E",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"7",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"6",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"7",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"6",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"7",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"E",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"6",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"E",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"7",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"9",    x"E",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"6",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"E",    x"9",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"7",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"E",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"6",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"E",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"7",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"D",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"A",    x"F",    x"F",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"D",    x"F",    x"F",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"D",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"6",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"D",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"F",    x"F",    x"D",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"F",    x"F",    x"A",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"7",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"D",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"A",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"6",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"A",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"7",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"A",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"E",    x"6",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"5",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"6",    x"6",    x"9",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"7",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"7",    x"E",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"A",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"7",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"4",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"2",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"4",    x"0",    x"0",    x"5",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"4",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"4",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"7",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"4",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"2",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"4",    x"0",    x"0",    x"5",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"4",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"4",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"7",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"4",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"2",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"4",    x"0",    x"0",    x"5",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"4",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"3",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"7",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"2",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"4",    x"0",    x"0",    x"5",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"4",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"7",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"2",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"4",    x"0",    x"0",    x"5",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"4",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"7",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"2",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"2",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"4",    x"0",    x"0",    x"5",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"4",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"2",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"7",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"2",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"2",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"4",    x"0",    x"0",    x"5",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"4",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"2",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"7",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"2",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"2",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"4",    x"0",    x"0",    x"5",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"4",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"2",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"7",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"2",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"2",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"4",    x"0",    x"0",    x"5",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"4",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"2",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"7",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"3",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"2",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"4",    x"0",    x"0",    x"5",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"4",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"3",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"7",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"3",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"2",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"4",    x"0",    x"0",    x"5",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"4",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"3",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"7",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"4",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"2",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"4",    x"0",    x"0",    x"5",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"4",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"7",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"4",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"2",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"4",    x"0",    x"0",    x"5",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"4",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"4",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"7",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"E",
        x"4",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"2",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"4",    x"0",    x"0",    x"5",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"4",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"4",
        x"E",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"7",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"6",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"2",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"4",    x"0",    x"0",    x"5",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"4",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"7",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"7",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"9",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"2",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"4",    x"0",    x"0",    x"5",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"4",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"8",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"7",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"2",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"4",    x"0",    x"0",    x"5",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"4",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"8",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"7",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"2",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"4",    x"0",    x"0",    x"5",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"4",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"7",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"1",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"2",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"4",    x"0",    x"0",    x"5",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"4",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"1",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"7",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"2",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"2",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"4",    x"0",    x"0",    x"5",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"4",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"2",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"7",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"2",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"4",    x"0",    x"0",    x"5",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"4",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"7",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"4",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"2",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"4",    x"0",    x"0",    x"5",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"4",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"4",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"7",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"5",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"2",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"4",    x"0",    x"0",    x"5",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"4",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"7",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"2",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"4",    x"0",    x"0",    x"5",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"4",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"7",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"1",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"2",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"4",    x"0",    x"0",    x"5",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"4",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"1",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"7",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"2",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"2",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"4",    x"0",    x"0",    x"5",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"4",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"2",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"7",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"4",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"2",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"4",    x"0",    x"0",    x"5",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"4",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"4",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"7",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"6",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"2",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"4",    x"0",    x"0",    x"5",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"4",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"6",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"7",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"2",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"4",    x"0",    x"0",    x"5",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"4",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"7",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"1",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"2",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"4",    x"0",    x"0",    x"5",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"4",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"1",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"7",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"2",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"4",    x"0",    x"0",    x"5",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"4",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"7",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"6",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"2",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"4",    x"0",    x"0",    x"5",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"4",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"7",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"5",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"2",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"4",    x"0",    x"0",    x"5",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"2",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"7",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"E",    x"F",
        x"E",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"D",    x"F",    x"F",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"B",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"2",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"4",    x"0",    x"0",    x"5",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"2",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"B",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"F",    x"F",    x"D",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"E",
        x"F",    x"E",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"2",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"2",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"4",    x"0",    x"0",    x"5",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"2",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"2",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"E",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"E",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"E",    x"F",    x"F",    x"E",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"A",    x"0",
        x"0",    x"0",    x"0",    x"6",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"6",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"6",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"A",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"E",    x"F",    x"F",    x"E",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"E",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"E",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"1",    x"0",
        x"0",    x"0",    x"0",    x"6",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"6",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"6",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"6",    x"8",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"3",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"6",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"6",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"6",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"6",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"6",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"6",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"6",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"6",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"6",    x"B",    x"A",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"6",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"6",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"6",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"6",    x"B",    x"B",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"6",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"6",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"6",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"6",    x"B",    x"B",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"6",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"6",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"6",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"6",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"6",    x"B",    x"B",    x"B",    x"A",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"1",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"6",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"6",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"6",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"6",    x"B",    x"B",    x"B",    x"B",    x"8",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"4",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"6",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"6",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"6",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"6",    x"B",    x"B",    x"B",    x"B",    x"B",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"6",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"6",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"6",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"6",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"6",    x"B",    x"B",    x"B",    x"B",    x"B",    x"A",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"1",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"6",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"6",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"6",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"6",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"8",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"5",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"6",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"6",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"6",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"6",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"6",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"6",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"6",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"6",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"9",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"2",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"6",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"6",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"6",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"6",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"6",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"6",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"6",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"6",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"6",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"A",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"1",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"6",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"6",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"6",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"6",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"5",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"6",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"6",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"6",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"6",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"6",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"6",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"6",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"6",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"4",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"6",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"6",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"6",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"6",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"6",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"6",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"6",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"6",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"9",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"2",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"6",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"6",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"6",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"6",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"6",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"6",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"6",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"6",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"6",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"1",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"6",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"6",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"6",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"6",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"6",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"6",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"6",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"6",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"6",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"A",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"1",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"6",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"6",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"6",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"6",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"5",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"6",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"6",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"6",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"6",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"A",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"1",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"6",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"6",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"6",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"6",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"8",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"5",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"6",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"6",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"6",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"6",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"6",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"6",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"6",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"6",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"8",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"5",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"6",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"6",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"6",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"6",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"6",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"6",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"6",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"6",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"9",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"5",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"6",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"6",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"6",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"6",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"E",    x"1",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"6",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"6",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"6",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"6",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"E",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"8",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"6",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"6",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"6",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"6",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"D",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"E",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"E",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"E",    x"E",    x"2",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"6",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"6",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"6",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"6",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"E",    x"E",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"E",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"E",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"B",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"7",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"7",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"7",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"7",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"7",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"7",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"7",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"7",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"D",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"E",    x"F",
        x"E",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"D",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"D",    x"9",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"9",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"6",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"6",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"6",    x"D",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"D",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"E",
        x"F",    x"E",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"9",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"6",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"6",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"9",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"9",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"9",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"6",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"6",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"8",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"9",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"6",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"6",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"9",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"9",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"6",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"6",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"9",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"6",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"6",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"4",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"9",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"9",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"6",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"6",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"8",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"9",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"6",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"6",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"6",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"9",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"6",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"6",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"9",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"6",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"6",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"9",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"6",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"6",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"4",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"9",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"6",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"6",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"9",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"6",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"6",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"6",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"9",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"6",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"6",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"9",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"9",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"6",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"6",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"9",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"6",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"6",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"5",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"9",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"6",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"6",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"9",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"9",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"6",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"6",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"9",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"6",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"6",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"5",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"8",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"9",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"6",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"6",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"8",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"9",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"9",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"6",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"6",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"8",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"9",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"6",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"6",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"4",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"8",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"9",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"6",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"6",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"8",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"9",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"9",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"6",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"6",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"8",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"9",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"6",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"6",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"4",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"8",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"9",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"6",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"6",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"9",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"9",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"6",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"6",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"8",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"9",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"6",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"6",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"6",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"9",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"6",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"6",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"9",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"9",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"6",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"6",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"9",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"9",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"6",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"6",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"8",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"9",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"6",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"6",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"4",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"9",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"6",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"6",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"9",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"6",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"6",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"9",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"9",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"6",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"6",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"6",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"E",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"9",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"6",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"6",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"4",    x"E",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"D",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"C",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"9",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"6",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"6",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"A",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"C",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"D",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"9",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"6",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"6",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"9",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"6",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"6",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"6",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"9",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"6",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"6",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"4",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"9",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"6",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"6",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"9",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"9",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"6",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"6",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"9",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"9",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"6",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"6",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"6",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"9",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"6",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"6",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"5",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"9",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"6",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"6",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"9",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"9",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"6",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"6",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"9",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"9",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"6",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"6",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"9",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"9",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"6",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"6",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"6",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"9",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"6",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"6",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"5",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"9",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"6",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"6",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"8",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"9",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"6",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"6",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"9",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"9",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"6",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"6",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"9",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"9",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"6",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"6",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"8",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"9",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"6",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"6",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"6",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"8",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"9",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"6",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"6",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"4",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"8",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"9",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"6",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"6",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"8",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"9",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"6",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"6",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"9",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"9",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"6",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"6",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"9",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"9",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"6",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"6",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"9",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"9",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"6",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"6",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"6",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"8",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"9",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"6",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"6",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"6",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"8",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"9",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"6",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"6",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"5",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"9",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"6",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"6",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"8",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"9",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"6",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"6",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"9",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"9",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"6",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"6",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"9",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"6",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"6",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"B",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"9",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"6",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"6",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"9",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"6",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"6",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"9",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"6",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"6",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"6",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"D",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"9",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"6",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"6",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"6",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"9",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"6",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"6",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"5",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"8",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"7",    x"A",    x"A",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"9",    x"A",    x"8",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"7",    x"A",    x"A",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"9",    x"A",    x"8",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"6",
        x"9",    x"9",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"9",    x"9",    x"8",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"8",    x"A",    x"9",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"A",    x"A",
        x"7",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"8",    x"9",    x"9",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"9",    x"9",    x"6",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"8",    x"9",    x"9",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"9",    x"9",    x"6",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"D",    x"F",
        x"D",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"B",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"9",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"5",    x"F",    x"F",    x"2",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"A",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"5",    x"F",    x"F",    x"2",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"A",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"5",
        x"F",    x"F",    x"2",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"C",    x"F",    x"A",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"A",    x"F",    x"C",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"2",    x"F",    x"F",
        x"5",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"A",    x"F",    x"C",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"2",    x"F",    x"F",    x"5",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"A",    x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"F",    x"F",    x"5",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"B",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"D",
        x"F",    x"D",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"5",    x"F",    x"F",    x"2",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"A",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"5",    x"F",    x"F",    x"2",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"A",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"5",
        x"F",    x"F",    x"2",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"C",    x"F",    x"A",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"A",    x"F",    x"C",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"2",    x"F",    x"F",
        x"5",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"A",    x"F",    x"C",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"2",    x"F",    x"F",    x"5",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"A",    x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"F",    x"F",    x"5",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"5",    x"F",    x"F",    x"2",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"A",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"5",    x"F",    x"F",    x"2",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"A",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"5",
        x"F",    x"F",    x"2",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"C",    x"F",    x"A",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"A",    x"F",    x"C",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"2",    x"F",    x"F",
        x"5",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"A",    x"F",    x"C",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"2",    x"F",    x"F",    x"5",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"A",    x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"F",    x"F",    x"5",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"5",    x"F",    x"F",    x"2",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"A",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"5",    x"F",    x"F",    x"2",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"A",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"5",
        x"F",    x"F",    x"2",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"C",    x"F",    x"A",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"A",    x"F",    x"C",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"2",    x"F",    x"F",
        x"5",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"A",    x"F",    x"C",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"2",    x"F",    x"F",    x"5",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"A",    x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"F",    x"F",    x"5",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"6",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"5",    x"F",    x"F",    x"2",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"A",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"5",    x"F",    x"F",    x"2",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"A",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"5",
        x"F",    x"F",    x"2",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"C",    x"F",    x"A",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"A",    x"F",    x"C",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"2",    x"F",    x"F",
        x"5",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"A",    x"F",    x"C",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"2",    x"F",    x"F",    x"5",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"A",    x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"F",    x"F",    x"5",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"6",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"6",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"5",    x"F",    x"F",    x"2",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"A",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"5",    x"F",    x"F",    x"2",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"A",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"5",
        x"F",    x"F",    x"2",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"C",    x"F",    x"A",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"A",    x"F",    x"C",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"2",    x"F",    x"F",
        x"5",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"A",    x"F",    x"C",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"2",    x"F",    x"F",    x"5",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"A",    x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"F",    x"F",    x"5",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"6",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"6",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"5",    x"F",    x"F",    x"2",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"A",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"5",    x"F",    x"F",    x"2",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"A",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"5",
        x"F",    x"F",    x"2",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"C",    x"F",    x"A",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"A",    x"F",    x"C",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"2",    x"F",    x"F",
        x"5",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"A",    x"F",    x"C",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"2",    x"F",    x"F",    x"5",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"A",    x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"F",    x"F",    x"5",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"6",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"6",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"5",    x"F",    x"F",    x"2",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"A",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"5",    x"F",    x"F",    x"2",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"A",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"5",
        x"F",    x"F",    x"2",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"C",    x"F",    x"A",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"A",    x"F",    x"C",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"2",    x"F",    x"F",
        x"5",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"A",    x"F",    x"C",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"2",    x"F",    x"F",    x"5",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"A",    x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"F",    x"F",    x"5",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"6",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"5",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"5",    x"F",    x"F",    x"2",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"A",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"5",    x"F",    x"F",    x"2",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"A",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"5",
        x"F",    x"F",    x"2",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"C",    x"F",    x"A",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"A",    x"F",    x"C",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"2",    x"F",    x"F",
        x"5",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"A",    x"F",    x"C",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"2",    x"F",    x"F",    x"5",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"A",    x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"F",    x"F",    x"5",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"6",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"5",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"5",    x"F",    x"F",    x"2",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"A",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"5",    x"F",    x"F",    x"2",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"A",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"5",
        x"F",    x"F",    x"2",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"C",    x"F",    x"A",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"A",    x"F",    x"C",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"2",    x"F",    x"F",
        x"5",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"A",    x"F",    x"C",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"2",    x"F",    x"F",    x"5",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"A",    x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"F",    x"F",    x"5",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"5",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"5",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"5",    x"F",    x"F",    x"2",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"A",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"5",    x"F",    x"F",    x"2",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"A",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"5",
        x"F",    x"F",    x"2",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"C",    x"F",    x"A",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"A",    x"F",    x"C",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"2",    x"F",    x"F",
        x"5",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"A",    x"F",    x"C",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"2",    x"F",    x"F",    x"5",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"A",    x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"F",    x"F",    x"5",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"5",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"5",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"5",    x"F",    x"F",    x"2",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"A",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"5",    x"F",    x"F",    x"2",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"A",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"5",
        x"F",    x"F",    x"2",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"C",    x"F",    x"A",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"A",    x"F",    x"C",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"2",    x"F",    x"F",
        x"5",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"A",    x"F",    x"C",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"2",    x"F",    x"F",    x"5",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"A",    x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"F",    x"F",    x"5",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"5",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"5",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"5",    x"F",    x"F",    x"2",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"A",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"5",    x"F",    x"F",    x"2",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"A",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"5",
        x"F",    x"F",    x"2",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"C",    x"F",    x"A",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"A",    x"F",    x"C",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"2",    x"F",    x"F",
        x"5",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"A",    x"F",    x"C",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"2",    x"F",    x"F",    x"5",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"A",    x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"F",    x"F",    x"5",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"5",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"5",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"5",    x"F",    x"F",    x"2",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"A",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"5",    x"F",    x"F",    x"2",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"A",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"5",
        x"F",    x"F",    x"2",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"C",    x"F",    x"A",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"A",    x"F",    x"C",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"2",    x"F",    x"F",
        x"5",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"A",    x"F",    x"C",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"2",    x"F",    x"F",    x"5",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"A",    x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"F",    x"F",    x"5",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"5",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"4",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"5",    x"F",    x"F",    x"2",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"A",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"5",    x"F",    x"F",    x"2",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"A",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"5",
        x"F",    x"F",    x"2",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"C",    x"F",    x"A",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"A",    x"F",    x"C",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"2",    x"F",    x"F",
        x"5",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"A",    x"F",    x"C",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"2",    x"F",    x"F",    x"5",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"A",    x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"F",    x"F",    x"5",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"4",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"5",    x"F",    x"F",    x"2",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"A",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"5",    x"F",    x"F",    x"2",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"A",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"5",
        x"F",    x"F",    x"2",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"C",    x"F",    x"A",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"A",    x"F",    x"C",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"2",    x"F",    x"F",
        x"5",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"A",    x"F",    x"C",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"2",    x"F",    x"F",    x"5",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"A",    x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"F",    x"F",    x"5",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"A",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"9",    x"F",    x"F",    x"7",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"D",    x"F",    x"C",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"9",    x"F",    x"F",    x"7",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"D",    x"F",    x"C",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"9",
        x"F",    x"F",    x"7",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"D",    x"F",    x"C",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"8",    x"F",
        x"F",    x"8",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"C",    x"F",    x"D",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",
        x"9",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"C",    x"F",    x"D",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"7",    x"F",    x"F",    x"9",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"C",    x"F",    x"D",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"7",    x"F",    x"F",    x"9",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"6",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"A",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"B",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"B",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"B",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"B",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"5",
        x"1",    x"1",    x"1",    x"1",    x"1",    x"1",    x"1",    x"1",
        x"1",    x"1",    x"1",    x"1",    x"1",    x"1",    x"1",    x"1",
        x"1",    x"5",    x"F",    x"F",    x"3",    x"1",    x"1",    x"1",
        x"1",    x"1",    x"1",    x"1",    x"1",    x"1",    x"1",    x"1",
        x"1",    x"1",    x"1",    x"1",    x"1",    x"1",    x"1",    x"1",
        x"1",    x"1",    x"1",    x"1",    x"1",    x"1",    x"1",    x"1",
        x"1",    x"1",    x"1",    x"1",    x"1",    x"C",    x"F",    x"A",
        x"1",    x"1",    x"1",    x"1",    x"1",    x"1",    x"1",    x"1",
        x"1",    x"1",    x"1",    x"1",    x"1",    x"1",    x"1",    x"1",
        x"1",    x"1",    x"1",    x"1",    x"1",    x"1",    x"1",    x"1",
        x"1",    x"1",    x"1",    x"1",    x"1",    x"1",    x"1",    x"1",
        x"5",    x"F",    x"F",    x"3",    x"1",    x"1",    x"1",    x"1",
        x"1",    x"1",    x"1",    x"1",    x"1",    x"1",    x"1",    x"1",
        x"1",    x"1",    x"1",    x"1",    x"1",    x"1",    x"1",    x"1",
        x"1",    x"1",    x"1",    x"1",    x"1",    x"1",    x"1",    x"1",
        x"1",    x"1",    x"1",    x"1",    x"C",    x"F",    x"A",    x"1",
        x"1",    x"1",    x"1",    x"1",    x"1",    x"1",    x"1",    x"1",
        x"1",    x"1",    x"1",    x"1",    x"1",    x"1",    x"1",    x"1",
        x"1",    x"1",    x"1",    x"1",    x"1",    x"1",    x"1",    x"1",
        x"1",    x"1",    x"1",    x"1",    x"1",    x"1",    x"1",    x"5",
        x"F",    x"F",    x"3",    x"1",    x"1",    x"1",    x"1",    x"1",
        x"1",    x"1",    x"1",    x"1",    x"1",    x"1",    x"1",    x"1",
        x"1",    x"1",    x"1",    x"1",    x"1",    x"1",    x"1",    x"1",
        x"1",    x"1",    x"1",    x"1",    x"1",    x"1",    x"1",    x"1",
        x"1",    x"1",    x"1",    x"C",    x"F",    x"A",    x"1",    x"1",
        x"1",    x"1",    x"1",    x"1",    x"1",    x"1",    x"1",    x"1",
        x"1",    x"1",    x"1",    x"1",    x"1",    x"1",    x"4",    x"F",
        x"F",    x"4",    x"1",    x"1",    x"1",    x"1",    x"1",    x"1",
        x"1",    x"1",    x"1",    x"1",    x"1",    x"1",    x"1",    x"1",
        x"1",    x"1",    x"A",    x"F",    x"C",    x"1",    x"1",    x"1",
        x"1",    x"1",    x"1",    x"1",    x"1",    x"1",    x"1",    x"1",
        x"1",    x"1",    x"1",    x"1",    x"1",    x"1",    x"1",    x"1",
        x"1",    x"1",    x"1",    x"1",    x"1",    x"1",    x"1",    x"1",
        x"1",    x"1",    x"1",    x"1",    x"1",    x"3",    x"F",    x"F",
        x"5",    x"1",    x"1",    x"1",    x"1",    x"1",    x"1",    x"1",
        x"1",    x"1",    x"1",    x"1",    x"1",    x"1",    x"1",    x"1",
        x"1",    x"1",    x"1",    x"1",    x"1",    x"1",    x"1",    x"1",
        x"1",    x"1",    x"1",    x"1",    x"1",    x"1",    x"1",    x"1",
        x"1",    x"A",    x"F",    x"C",    x"1",    x"1",    x"1",    x"1",
        x"1",    x"1",    x"1",    x"1",    x"1",    x"1",    x"1",    x"1",
        x"1",    x"1",    x"1",    x"1",    x"1",    x"1",    x"1",    x"1",
        x"1",    x"1",    x"1",    x"1",    x"1",    x"1",    x"1",    x"1",
        x"1",    x"1",    x"1",    x"1",    x"3",    x"F",    x"F",    x"5",
        x"1",    x"1",    x"1",    x"1",    x"1",    x"1",    x"1",    x"1",
        x"1",    x"1",    x"1",    x"1",    x"1",    x"1",    x"1",    x"1",
        x"1",    x"1",    x"1",    x"1",    x"1",    x"1",    x"1",    x"1",
        x"1",    x"1",    x"1",    x"1",    x"1",    x"1",    x"1",    x"1",
        x"A",    x"F",    x"C",    x"1",    x"1",    x"1",    x"1",    x"1",
        x"1",    x"1",    x"1",    x"1",    x"1",    x"1",    x"1",    x"1",
        x"1",    x"1",    x"1",    x"1",    x"1",    x"1",    x"1",    x"1",
        x"1",    x"1",    x"1",    x"1",    x"1",    x"1",    x"1",    x"1",
        x"1",    x"1",    x"1",    x"3",    x"F",    x"F",    x"5",    x"1",
        x"1",    x"1",    x"1",    x"1",    x"1",    x"1",    x"1",    x"1",
        x"1",    x"1",    x"1",    x"1",    x"1",    x"1",    x"1",    x"1",
        x"5",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"5",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"5",    x"F",    x"F",    x"2",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"A",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"5",    x"F",    x"F",    x"2",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"A",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"5",
        x"F",    x"F",    x"2",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"C",    x"F",    x"A",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"A",    x"F",    x"C",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"2",    x"F",    x"F",
        x"5",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"A",    x"F",    x"C",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"2",    x"F",    x"F",    x"5",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"A",    x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"F",    x"F",    x"5",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"5",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"5",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"5",    x"F",    x"F",    x"2",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"A",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"5",    x"F",    x"F",    x"2",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"A",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"5",
        x"F",    x"F",    x"2",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"C",    x"F",    x"A",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"A",    x"F",    x"C",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"2",    x"F",    x"F",
        x"5",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"A",    x"F",    x"C",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"2",    x"F",    x"F",    x"5",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"A",    x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"F",    x"F",    x"5",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"5",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"5",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"5",    x"F",    x"F",    x"2",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"A",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"5",    x"F",    x"F",    x"2",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"A",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"5",
        x"F",    x"F",    x"2",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"C",    x"F",    x"A",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"A",    x"F",    x"C",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"2",    x"F",    x"F",
        x"5",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"A",    x"F",    x"C",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"2",    x"F",    x"F",    x"5",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"A",    x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"F",    x"F",    x"5",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"5",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"5",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"5",    x"F",    x"F",    x"2",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"A",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"5",    x"F",    x"F",    x"2",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"A",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"5",
        x"F",    x"F",    x"2",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"C",    x"F",    x"A",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"A",    x"F",    x"C",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"2",    x"F",    x"F",
        x"5",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"A",    x"F",    x"C",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"2",    x"F",    x"F",    x"5",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"A",    x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"F",    x"F",    x"5",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"5",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"5",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"5",    x"F",    x"F",    x"2",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"A",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"5",    x"F",    x"F",    x"2",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"A",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"5",
        x"F",    x"F",    x"2",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"C",    x"F",    x"A",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"A",    x"F",    x"C",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"2",    x"F",    x"F",
        x"5",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"A",    x"F",    x"C",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"2",    x"F",    x"F",    x"5",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"A",    x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"F",    x"F",    x"5",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"5",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"5",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"5",    x"F",    x"F",    x"2",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"A",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"5",    x"F",    x"F",    x"2",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"A",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"5",
        x"F",    x"F",    x"2",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"C",    x"F",    x"A",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"A",    x"F",    x"C",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"2",    x"F",    x"F",
        x"5",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"A",    x"F",    x"C",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"2",    x"F",    x"F",    x"5",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"A",    x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"F",    x"F",    x"5",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"6",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"6",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"5",    x"F",    x"F",    x"2",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"A",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"5",    x"F",    x"F",    x"2",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"A",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"5",
        x"F",    x"F",    x"2",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"C",    x"F",    x"A",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"A",    x"F",    x"C",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"2",    x"F",    x"F",
        x"5",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"A",    x"F",    x"C",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"2",    x"F",    x"F",    x"5",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"A",    x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"F",    x"F",    x"5",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"6",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"6",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"5",    x"F",    x"F",    x"2",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"A",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"5",    x"F",    x"F",    x"2",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"A",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"5",
        x"F",    x"F",    x"2",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"C",    x"F",    x"A",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"A",    x"F",    x"C",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"2",    x"F",    x"F",
        x"5",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"A",    x"F",    x"C",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"2",    x"F",    x"F",    x"5",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"A",    x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"F",    x"F",    x"5",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"6",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"6",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"5",    x"F",    x"F",    x"2",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"A",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"5",    x"F",    x"F",    x"2",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"A",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"5",
        x"F",    x"F",    x"2",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"C",    x"F",    x"A",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"A",    x"F",    x"C",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"2",    x"F",    x"F",
        x"5",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"A",    x"F",    x"C",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"2",    x"F",    x"F",    x"5",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"A",    x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"F",    x"F",    x"5",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"6",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"6",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"5",    x"F",    x"F",    x"2",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"A",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"5",    x"F",    x"F",    x"2",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"A",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"5",
        x"F",    x"F",    x"2",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"C",    x"F",    x"A",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"A",    x"F",    x"C",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"2",    x"F",    x"F",
        x"5",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"A",    x"F",    x"C",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"2",    x"F",    x"F",    x"5",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"A",    x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"F",    x"F",    x"5",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"6",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"5",    x"F",    x"F",    x"2",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"A",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"5",    x"F",    x"F",    x"2",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"A",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"5",
        x"F",    x"F",    x"2",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"C",    x"F",    x"A",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"A",    x"F",    x"C",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"2",    x"F",    x"F",
        x"5",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"A",    x"F",    x"C",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"2",    x"F",    x"F",    x"5",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"A",    x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"F",    x"F",    x"5",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"5",    x"F",    x"F",    x"2",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"A",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"5",    x"F",    x"F",    x"2",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"A",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"5",
        x"F",    x"F",    x"2",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"C",    x"F",    x"A",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"A",    x"F",    x"C",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"2",    x"F",    x"F",
        x"5",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"A",    x"F",    x"C",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"2",    x"F",    x"F",    x"5",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"A",    x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"F",    x"F",    x"5",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"5",    x"F",    x"F",    x"2",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"A",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"5",    x"F",    x"F",    x"2",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"A",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"5",
        x"F",    x"F",    x"2",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"C",    x"F",    x"A",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"A",    x"F",    x"C",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"2",    x"F",    x"F",
        x"5",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"A",    x"F",    x"C",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"2",    x"F",    x"F",    x"5",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"A",    x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"F",    x"F",    x"5",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"D",    x"F",
        x"D",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"B",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"5",    x"F",    x"F",    x"2",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"A",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"5",    x"F",    x"F",    x"2",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"A",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"5",
        x"F",    x"F",    x"2",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"C",    x"F",    x"A",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"A",    x"F",    x"C",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"2",    x"F",    x"F",
        x"5",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"A",    x"F",    x"C",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"2",    x"F",    x"F",    x"5",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"A",    x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"F",    x"F",    x"5",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"B",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"D",
        x"F",    x"D",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"5",    x"F",    x"F",    x"2",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"A",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"5",    x"F",    x"F",    x"2",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"A",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"5",
        x"F",    x"F",    x"2",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"C",    x"F",    x"A",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"A",    x"F",    x"C",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"2",    x"F",    x"F",
        x"5",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"A",    x"F",    x"C",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"2",    x"F",    x"F",    x"5",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"A",    x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"F",    x"F",    x"5",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"1",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"1",    x"5",    x"5",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"1",    x"3",    x"4",    x"5",    x"6",
        x"7",    x"8",    x"9",    x"8",    x"7",    x"6",    x"5",    x"4",
        x"2",    x"1",    x"0",    x"0",    x"1",    x"6",    x"7",    x"7",
        x"6",    x"7",    x"9",    x"9",    x"8",    x"7",    x"6",    x"5",
        x"3",    x"2",    x"1",    x"0",    x"0",    x"2",    x"3",    x"4",
        x"5",    x"6",    x"8",    x"9",    x"9",    x"8",    x"7",    x"6",
        x"4",    x"3",    x"2",    x"1",    x"0",    x"1",    x"2",    x"3",
        x"5",    x"8",    x"9",    x"8",    x"9",    x"9",    x"8",    x"7",
        x"5",    x"4",    x"3",    x"2",    x"1",    x"0",    x"1",    x"2",
        x"3",    x"4",    x"6",    x"7",    x"8",    x"9",    x"9",    x"8",
        x"6",    x"5",    x"4",    x"3",    x"4",    x"5",    x"8",    x"8",
        x"5",    x"2",    x"0",    x"3",    x"8",    x"B",    x"9",    x"4",
        x"1",    x"1",    x"4",    x"7",    x"9",    x"7",    x"4",    x"1",
        x"1",    x"4",    x"7",    x"9",    x"6",    x"3",    x"0",    x"2",
        x"5",    x"8",    x"8",    x"5",    x"2",    x"0",    x"3",    x"6",
        x"9",    x"7",    x"4",    x"1",    x"1",    x"4",    x"7",    x"A",
        x"9",    x"7",    x"1",    x"1",    x"4",    x"7",    x"9",    x"6",
        x"3",    x"0",    x"2",    x"5",    x"8",    x"8",    x"5",    x"2",
        x"0",    x"3",    x"6",    x"9",    x"7",    x"4",    x"1",    x"5",
        x"8",    x"8",    x"6",    x"3",    x"5",    x"8",    x"8",    x"6",
        x"3",    x"5",    x"8",    x"A",    x"9",    x"5",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"A",    x"A",    x"8",    x"3",    x"6",    x"9",
        x"8",    x"5",    x"3",    x"6",    x"9",    x"8",    x"5",    x"4",
        x"6",    x"9",    x"7",    x"5",    x"4",    x"6",    x"9",    x"7",
        x"5",    x"2",    x"8",    x"5",    x"0",    x"6",    x"7",    x"1",
        x"4",    x"9",    x"3",    x"2",    x"8",    x"6",    x"5",    x"9",
        x"8",    x"1",    x"4",    x"A",    x"4",    x"2",    x"8",    x"6",
        x"0",    x"5",    x"8",    x"2",    x"3",    x"9",    x"4",    x"1",
        x"7",    x"6",    x"0",    x"5",    x"8",    x"2",    x"3",    x"9",
        x"4",    x"1",    x"7",    x"6",    x"0",    x"5",    x"8",    x"2",
        x"3",    x"B",    x"7",    x"5",    x"7",    x"6",    x"0",    x"5",
        x"8",    x"2",    x"3",    x"9",    x"4",    x"1",    x"7",    x"6",
        x"0",    x"5",    x"8",    x"2",    x"3",    x"9",    x"4",    x"1",
        x"7",    x"6",    x"0",    x"5",    x"8",    x"2",    x"3",    x"9",
        x"4",    x"6",    x"0",    x"8",    x"4",    x"7",    x"A",    x"2",
        x"8",    x"3",    x"4",    x"7",    x"0",    x"8",    x"3",    x"4",
        x"7",    x"1",    x"9",    x"2",    x"5",    x"6",    x"1",    x"9",
        x"2",    x"5",    x"6",    x"1",    x"9",    x"2",    x"5",    x"6",
        x"2",    x"9",    x"1",    x"6",    x"5",    x"2",    x"9",    x"1",
        x"8",    x"8",    x"6",    x"9",    x"1",    x"6",    x"5",    x"3",
        x"9",    x"0",    x"7",    x"4",    x"3",    x"8",    x"0",    x"7",
        x"4",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"5",    x"5",    x"1",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"1",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"4",    x"6",    x"8",    x"9",
        x"B",    x"D",    x"E",    x"D",    x"B",    x"9",    x"7",    x"6",
        x"4",    x"2",    x"0",    x"1",    x"2",    x"4",    x"6",    x"8",
        x"A",    x"B",    x"D",    x"E",    x"C",    x"B",    x"9",    x"7",
        x"5",    x"3",    x"2",    x"0",    x"1",    x"3",    x"4",    x"6",
        x"8",    x"A",    x"C",    x"D",    x"E",    x"C",    x"A",    x"9",
        x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",    x"5",
        x"7",    x"8",    x"A",    x"C",    x"E",    x"E",    x"C",    x"A",
        x"8",    x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",
        x"5",    x"7",    x"9",    x"A",    x"C",    x"E",    x"D",    x"C",
        x"A",    x"8",    x"6",    x"5",    x"6",    x"8",    x"C",    x"C",
        x"8",    x"4",    x"0",    x"4",    x"9",    x"D",    x"B",    x"7",
        x"2",    x"1",    x"6",    x"A",    x"E",    x"A",    x"6",    x"1",
        x"2",    x"7",    x"B",    x"D",    x"9",    x"5",    x"0",    x"3",
        x"8",    x"C",    x"C",    x"8",    x"3",    x"0",    x"5",    x"9",
        x"D",    x"B",    x"7",    x"2",    x"1",    x"6",    x"A",    x"E",
        x"A",    x"6",    x"1",    x"2",    x"7",    x"B",    x"D",    x"9",
        x"4",    x"0",    x"4",    x"8",    x"D",    x"C",    x"8",    x"3",
        x"0",    x"5",    x"9",    x"E",    x"B",    x"6",    x"0",    x"5",
        x"B",    x"C",    x"6",    x"0",    x"5",    x"B",    x"C",    x"6",
        x"0",    x"5",    x"B",    x"C",    x"6",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",
        x"A",    x"4",    x"1",    x"7",    x"D",    x"A",    x"4",    x"1",
        x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",    x"A",
        x"4",    x"2",    x"C",    x"8",    x"0",    x"9",    x"B",    x"2",
        x"6",    x"E",    x"5",    x"3",    x"C",    x"8",    x"0",    x"9",
        x"B",    x"2",    x"6",    x"F",    x"6",    x"3",    x"C",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"2",    x"B",    x"9",    x"0",    x"8",    x"C",    x"3",
        x"5",    x"E",    x"6",    x"2",    x"B",    x"9",    x"0",    x"8",
        x"C",    x"3",    x"5",    x"E",    x"6",    x"2",    x"B",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"9",    x"0",    x"C",    x"5",    x"6",    x"B",    x"0",
        x"C",    x"5",    x"6",    x"B",    x"1",    x"D",    x"4",    x"7",
        x"A",    x"1",    x"D",    x"4",    x"7",    x"A",    x"2",    x"E",
        x"3",    x"8",    x"9",    x"2",    x"E",    x"3",    x"8",    x"9",
        x"3",    x"E",    x"2",    x"9",    x"8",    x"3",    x"E",    x"2",
        x"9",    x"8",    x"4",    x"D",    x"1",    x"A",    x"7",    x"4",
        x"D",    x"1",    x"A",    x"7",    x"4",    x"C",    x"0",    x"B",
        x"6",    x"1",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"4",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"4",    x"6",    x"8",    x"9",
        x"B",    x"D",    x"E",    x"D",    x"B",    x"9",    x"7",    x"6",
        x"4",    x"2",    x"0",    x"1",    x"2",    x"4",    x"6",    x"8",
        x"A",    x"B",    x"D",    x"E",    x"C",    x"B",    x"9",    x"7",
        x"5",    x"3",    x"2",    x"0",    x"1",    x"3",    x"4",    x"6",
        x"8",    x"A",    x"C",    x"D",    x"E",    x"C",    x"A",    x"9",
        x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",    x"5",
        x"7",    x"8",    x"A",    x"C",    x"E",    x"E",    x"C",    x"A",
        x"8",    x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",
        x"5",    x"7",    x"9",    x"A",    x"C",    x"E",    x"D",    x"C",
        x"A",    x"8",    x"6",    x"5",    x"6",    x"8",    x"C",    x"C",
        x"8",    x"4",    x"0",    x"4",    x"9",    x"D",    x"B",    x"7",
        x"2",    x"1",    x"6",    x"A",    x"E",    x"A",    x"6",    x"1",
        x"2",    x"7",    x"B",    x"D",    x"9",    x"5",    x"0",    x"3",
        x"8",    x"C",    x"C",    x"8",    x"3",    x"0",    x"5",    x"9",
        x"D",    x"B",    x"7",    x"2",    x"1",    x"6",    x"A",    x"E",
        x"A",    x"6",    x"1",    x"2",    x"7",    x"B",    x"D",    x"9",
        x"4",    x"0",    x"4",    x"8",    x"D",    x"C",    x"8",    x"3",
        x"0",    x"5",    x"9",    x"E",    x"B",    x"6",    x"0",    x"5",
        x"B",    x"C",    x"6",    x"0",    x"5",    x"B",    x"C",    x"6",
        x"0",    x"5",    x"B",    x"C",    x"6",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",
        x"A",    x"4",    x"1",    x"7",    x"D",    x"A",    x"4",    x"1",
        x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",    x"A",
        x"4",    x"2",    x"C",    x"8",    x"0",    x"9",    x"B",    x"2",
        x"6",    x"E",    x"5",    x"3",    x"C",    x"8",    x"0",    x"9",
        x"B",    x"2",    x"6",    x"F",    x"6",    x"3",    x"C",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"2",    x"B",    x"9",    x"0",    x"8",    x"C",    x"3",
        x"5",    x"E",    x"6",    x"2",    x"B",    x"9",    x"0",    x"8",
        x"C",    x"3",    x"5",    x"E",    x"6",    x"2",    x"B",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"9",    x"0",    x"C",    x"5",    x"6",    x"B",    x"0",
        x"C",    x"5",    x"6",    x"B",    x"1",    x"D",    x"4",    x"7",
        x"A",    x"1",    x"D",    x"4",    x"7",    x"A",    x"2",    x"E",
        x"3",    x"8",    x"9",    x"2",    x"E",    x"3",    x"8",    x"9",
        x"3",    x"E",    x"2",    x"9",    x"8",    x"3",    x"E",    x"2",
        x"9",    x"8",    x"4",    x"D",    x"1",    x"A",    x"7",    x"4",
        x"D",    x"1",    x"A",    x"7",    x"4",    x"C",    x"0",    x"B",
        x"6",    x"1",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"4",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"4",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"4",    x"6",    x"8",    x"9",
        x"B",    x"D",    x"E",    x"D",    x"B",    x"9",    x"7",    x"6",
        x"4",    x"2",    x"0",    x"1",    x"2",    x"4",    x"6",    x"8",
        x"A",    x"B",    x"D",    x"E",    x"C",    x"B",    x"9",    x"7",
        x"5",    x"3",    x"2",    x"0",    x"1",    x"3",    x"4",    x"6",
        x"8",    x"A",    x"C",    x"D",    x"E",    x"C",    x"A",    x"9",
        x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",    x"5",
        x"7",    x"8",    x"A",    x"C",    x"E",    x"E",    x"C",    x"A",
        x"8",    x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",
        x"5",    x"7",    x"9",    x"A",    x"C",    x"E",    x"D",    x"C",
        x"A",    x"8",    x"6",    x"5",    x"6",    x"8",    x"C",    x"C",
        x"8",    x"4",    x"0",    x"4",    x"9",    x"D",    x"B",    x"7",
        x"2",    x"1",    x"6",    x"A",    x"E",    x"A",    x"6",    x"1",
        x"2",    x"7",    x"B",    x"D",    x"9",    x"5",    x"0",    x"3",
        x"8",    x"C",    x"C",    x"8",    x"3",    x"0",    x"5",    x"9",
        x"D",    x"B",    x"7",    x"2",    x"1",    x"6",    x"A",    x"E",
        x"A",    x"6",    x"1",    x"2",    x"7",    x"B",    x"D",    x"9",
        x"4",    x"0",    x"4",    x"8",    x"D",    x"C",    x"8",    x"3",
        x"0",    x"5",    x"9",    x"E",    x"B",    x"6",    x"0",    x"5",
        x"B",    x"C",    x"6",    x"0",    x"5",    x"B",    x"C",    x"6",
        x"0",    x"5",    x"B",    x"C",    x"6",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",
        x"A",    x"4",    x"1",    x"7",    x"D",    x"A",    x"4",    x"1",
        x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",    x"A",
        x"4",    x"2",    x"C",    x"8",    x"0",    x"9",    x"B",    x"2",
        x"6",    x"E",    x"5",    x"3",    x"C",    x"8",    x"0",    x"9",
        x"B",    x"2",    x"6",    x"F",    x"6",    x"3",    x"C",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"2",    x"B",    x"9",    x"0",    x"8",    x"C",    x"3",
        x"5",    x"E",    x"6",    x"2",    x"B",    x"9",    x"0",    x"8",
        x"C",    x"3",    x"5",    x"E",    x"6",    x"2",    x"B",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"9",    x"0",    x"C",    x"5",    x"6",    x"B",    x"0",
        x"C",    x"5",    x"6",    x"B",    x"1",    x"D",    x"4",    x"7",
        x"A",    x"1",    x"D",    x"4",    x"7",    x"A",    x"2",    x"E",
        x"3",    x"8",    x"9",    x"2",    x"E",    x"3",    x"8",    x"9",
        x"3",    x"E",    x"2",    x"9",    x"8",    x"3",    x"E",    x"2",
        x"9",    x"8",    x"4",    x"D",    x"1",    x"A",    x"7",    x"4",
        x"D",    x"1",    x"A",    x"7",    x"4",    x"C",    x"0",    x"B",
        x"6",    x"1",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"4",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"5",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"4",    x"6",    x"8",    x"9",
        x"B",    x"D",    x"E",    x"D",    x"B",    x"9",    x"7",    x"6",
        x"4",    x"2",    x"0",    x"1",    x"2",    x"4",    x"6",    x"8",
        x"A",    x"B",    x"D",    x"E",    x"C",    x"B",    x"9",    x"7",
        x"5",    x"3",    x"2",    x"0",    x"1",    x"3",    x"4",    x"6",
        x"8",    x"A",    x"C",    x"D",    x"E",    x"C",    x"A",    x"9",
        x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",    x"5",
        x"7",    x"8",    x"A",    x"C",    x"E",    x"E",    x"C",    x"A",
        x"8",    x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",
        x"5",    x"7",    x"9",    x"A",    x"C",    x"E",    x"D",    x"C",
        x"A",    x"8",    x"6",    x"5",    x"6",    x"8",    x"C",    x"C",
        x"8",    x"4",    x"0",    x"4",    x"9",    x"D",    x"B",    x"7",
        x"2",    x"1",    x"6",    x"A",    x"E",    x"A",    x"6",    x"1",
        x"2",    x"7",    x"B",    x"D",    x"9",    x"5",    x"0",    x"3",
        x"8",    x"C",    x"C",    x"8",    x"3",    x"0",    x"5",    x"9",
        x"D",    x"B",    x"7",    x"2",    x"1",    x"6",    x"A",    x"E",
        x"A",    x"6",    x"1",    x"2",    x"7",    x"B",    x"D",    x"9",
        x"4",    x"0",    x"4",    x"8",    x"D",    x"C",    x"8",    x"3",
        x"0",    x"5",    x"9",    x"E",    x"B",    x"6",    x"0",    x"5",
        x"B",    x"C",    x"6",    x"0",    x"5",    x"B",    x"C",    x"6",
        x"0",    x"5",    x"B",    x"C",    x"6",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",
        x"A",    x"4",    x"1",    x"7",    x"D",    x"A",    x"4",    x"1",
        x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",    x"A",
        x"4",    x"2",    x"C",    x"8",    x"0",    x"9",    x"B",    x"2",
        x"6",    x"E",    x"5",    x"3",    x"C",    x"8",    x"0",    x"9",
        x"B",    x"2",    x"6",    x"F",    x"6",    x"3",    x"C",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"2",    x"B",    x"9",    x"0",    x"8",    x"C",    x"3",
        x"5",    x"E",    x"6",    x"2",    x"B",    x"9",    x"0",    x"8",
        x"C",    x"3",    x"5",    x"E",    x"6",    x"2",    x"B",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"9",    x"0",    x"C",    x"5",    x"6",    x"B",    x"0",
        x"C",    x"5",    x"6",    x"B",    x"1",    x"D",    x"4",    x"7",
        x"A",    x"1",    x"D",    x"4",    x"7",    x"A",    x"2",    x"E",
        x"3",    x"8",    x"9",    x"2",    x"E",    x"3",    x"8",    x"9",
        x"3",    x"E",    x"2",    x"9",    x"8",    x"3",    x"E",    x"2",
        x"9",    x"8",    x"4",    x"D",    x"1",    x"A",    x"7",    x"4",
        x"D",    x"1",    x"A",    x"7",    x"4",    x"C",    x"0",    x"B",
        x"6",    x"1",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"5",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"6",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"4",    x"6",    x"8",    x"9",
        x"B",    x"D",    x"E",    x"D",    x"B",    x"9",    x"7",    x"6",
        x"4",    x"2",    x"0",    x"1",    x"2",    x"4",    x"6",    x"8",
        x"A",    x"B",    x"D",    x"E",    x"C",    x"B",    x"9",    x"7",
        x"5",    x"3",    x"2",    x"0",    x"1",    x"3",    x"4",    x"6",
        x"8",    x"A",    x"C",    x"D",    x"E",    x"C",    x"A",    x"9",
        x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",    x"5",
        x"7",    x"8",    x"A",    x"C",    x"E",    x"E",    x"C",    x"A",
        x"8",    x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",
        x"5",    x"7",    x"9",    x"A",    x"C",    x"E",    x"D",    x"C",
        x"A",    x"8",    x"6",    x"5",    x"6",    x"8",    x"C",    x"C",
        x"8",    x"4",    x"0",    x"4",    x"9",    x"D",    x"B",    x"7",
        x"2",    x"1",    x"6",    x"A",    x"E",    x"A",    x"6",    x"1",
        x"2",    x"7",    x"B",    x"D",    x"9",    x"5",    x"0",    x"3",
        x"8",    x"C",    x"C",    x"8",    x"3",    x"0",    x"5",    x"9",
        x"D",    x"B",    x"7",    x"2",    x"1",    x"6",    x"A",    x"E",
        x"A",    x"6",    x"1",    x"2",    x"7",    x"B",    x"D",    x"9",
        x"4",    x"0",    x"4",    x"8",    x"D",    x"C",    x"8",    x"3",
        x"0",    x"5",    x"9",    x"E",    x"B",    x"6",    x"0",    x"5",
        x"B",    x"C",    x"6",    x"0",    x"5",    x"B",    x"C",    x"6",
        x"0",    x"5",    x"B",    x"C",    x"6",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",
        x"A",    x"4",    x"1",    x"7",    x"D",    x"A",    x"4",    x"1",
        x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",    x"A",
        x"4",    x"2",    x"C",    x"8",    x"0",    x"9",    x"B",    x"2",
        x"6",    x"E",    x"5",    x"3",    x"C",    x"8",    x"0",    x"9",
        x"B",    x"2",    x"6",    x"F",    x"6",    x"3",    x"C",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"2",    x"B",    x"9",    x"0",    x"8",    x"C",    x"3",
        x"5",    x"E",    x"6",    x"2",    x"B",    x"9",    x"0",    x"8",
        x"C",    x"3",    x"5",    x"E",    x"6",    x"2",    x"B",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"9",    x"0",    x"C",    x"5",    x"6",    x"B",    x"0",
        x"C",    x"5",    x"6",    x"B",    x"1",    x"D",    x"4",    x"7",
        x"A",    x"1",    x"D",    x"4",    x"7",    x"A",    x"2",    x"E",
        x"3",    x"8",    x"9",    x"2",    x"E",    x"3",    x"8",    x"9",
        x"3",    x"E",    x"2",    x"9",    x"8",    x"3",    x"E",    x"2",
        x"9",    x"8",    x"4",    x"D",    x"1",    x"A",    x"7",    x"4",
        x"D",    x"1",    x"A",    x"7",    x"4",    x"C",    x"0",    x"B",
        x"6",    x"1",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"4",    x"6",    x"8",    x"9",
        x"B",    x"D",    x"E",    x"D",    x"B",    x"9",    x"7",    x"6",
        x"4",    x"2",    x"0",    x"1",    x"2",    x"4",    x"6",    x"8",
        x"A",    x"B",    x"D",    x"E",    x"C",    x"B",    x"9",    x"7",
        x"5",    x"3",    x"2",    x"0",    x"1",    x"3",    x"4",    x"6",
        x"8",    x"A",    x"C",    x"D",    x"E",    x"C",    x"A",    x"9",
        x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",    x"5",
        x"7",    x"8",    x"A",    x"C",    x"E",    x"E",    x"C",    x"A",
        x"8",    x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",
        x"5",    x"7",    x"9",    x"A",    x"C",    x"E",    x"D",    x"C",
        x"A",    x"8",    x"6",    x"5",    x"6",    x"8",    x"C",    x"C",
        x"8",    x"4",    x"0",    x"4",    x"9",    x"D",    x"B",    x"7",
        x"2",    x"1",    x"6",    x"A",    x"E",    x"A",    x"6",    x"1",
        x"2",    x"7",    x"B",    x"D",    x"9",    x"5",    x"0",    x"3",
        x"8",    x"C",    x"C",    x"8",    x"3",    x"0",    x"5",    x"9",
        x"D",    x"B",    x"7",    x"2",    x"1",    x"6",    x"A",    x"E",
        x"A",    x"6",    x"1",    x"2",    x"7",    x"B",    x"D",    x"9",
        x"4",    x"0",    x"4",    x"8",    x"D",    x"C",    x"8",    x"3",
        x"0",    x"5",    x"9",    x"E",    x"B",    x"6",    x"0",    x"5",
        x"B",    x"C",    x"6",    x"0",    x"5",    x"B",    x"C",    x"6",
        x"0",    x"5",    x"B",    x"C",    x"6",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",
        x"A",    x"4",    x"1",    x"7",    x"D",    x"A",    x"4",    x"1",
        x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",    x"A",
        x"4",    x"2",    x"C",    x"8",    x"0",    x"9",    x"B",    x"2",
        x"6",    x"E",    x"5",    x"3",    x"C",    x"8",    x"0",    x"9",
        x"B",    x"2",    x"6",    x"F",    x"6",    x"3",    x"C",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"2",    x"B",    x"9",    x"0",    x"8",    x"C",    x"3",
        x"5",    x"E",    x"6",    x"2",    x"B",    x"9",    x"0",    x"8",
        x"C",    x"3",    x"5",    x"E",    x"6",    x"2",    x"B",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"9",    x"0",    x"C",    x"5",    x"6",    x"B",    x"0",
        x"C",    x"5",    x"6",    x"B",    x"1",    x"D",    x"4",    x"7",
        x"A",    x"1",    x"D",    x"4",    x"7",    x"A",    x"2",    x"E",
        x"3",    x"8",    x"9",    x"2",    x"E",    x"3",    x"8",    x"9",
        x"3",    x"E",    x"2",    x"9",    x"8",    x"3",    x"E",    x"2",
        x"9",    x"8",    x"4",    x"D",    x"1",    x"A",    x"7",    x"4",
        x"D",    x"1",    x"A",    x"7",    x"4",    x"C",    x"0",    x"B",
        x"6",    x"1",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"4",    x"6",    x"8",    x"9",
        x"B",    x"D",    x"E",    x"D",    x"B",    x"9",    x"7",    x"6",
        x"4",    x"2",    x"0",    x"1",    x"2",    x"4",    x"6",    x"8",
        x"A",    x"B",    x"D",    x"E",    x"C",    x"B",    x"9",    x"7",
        x"5",    x"3",    x"2",    x"0",    x"1",    x"3",    x"4",    x"6",
        x"8",    x"A",    x"C",    x"D",    x"E",    x"C",    x"A",    x"9",
        x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",    x"5",
        x"7",    x"8",    x"A",    x"C",    x"E",    x"E",    x"C",    x"A",
        x"8",    x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",
        x"5",    x"7",    x"9",    x"A",    x"C",    x"E",    x"D",    x"C",
        x"A",    x"8",    x"6",    x"5",    x"6",    x"8",    x"C",    x"C",
        x"8",    x"4",    x"0",    x"4",    x"9",    x"D",    x"B",    x"7",
        x"2",    x"1",    x"6",    x"A",    x"E",    x"A",    x"6",    x"1",
        x"2",    x"7",    x"B",    x"D",    x"9",    x"5",    x"0",    x"3",
        x"8",    x"C",    x"C",    x"8",    x"3",    x"0",    x"5",    x"9",
        x"D",    x"B",    x"7",    x"2",    x"1",    x"6",    x"A",    x"E",
        x"A",    x"6",    x"1",    x"2",    x"7",    x"B",    x"D",    x"9",
        x"4",    x"0",    x"4",    x"8",    x"D",    x"C",    x"8",    x"3",
        x"0",    x"5",    x"9",    x"E",    x"B",    x"6",    x"0",    x"5",
        x"B",    x"C",    x"6",    x"0",    x"5",    x"B",    x"C",    x"6",
        x"0",    x"5",    x"B",    x"C",    x"6",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",
        x"A",    x"4",    x"1",    x"7",    x"D",    x"A",    x"4",    x"1",
        x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",    x"A",
        x"4",    x"2",    x"C",    x"8",    x"0",    x"9",    x"B",    x"2",
        x"6",    x"E",    x"5",    x"3",    x"C",    x"8",    x"0",    x"9",
        x"B",    x"2",    x"6",    x"F",    x"6",    x"3",    x"C",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"2",    x"B",    x"9",    x"0",    x"8",    x"C",    x"3",
        x"5",    x"E",    x"6",    x"2",    x"B",    x"9",    x"0",    x"8",
        x"C",    x"3",    x"5",    x"E",    x"6",    x"2",    x"B",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"9",    x"0",    x"C",    x"5",    x"6",    x"B",    x"0",
        x"C",    x"5",    x"6",    x"B",    x"1",    x"D",    x"4",    x"7",
        x"A",    x"1",    x"D",    x"4",    x"7",    x"A",    x"2",    x"E",
        x"3",    x"8",    x"9",    x"2",    x"E",    x"3",    x"8",    x"9",
        x"3",    x"E",    x"2",    x"9",    x"8",    x"3",    x"E",    x"2",
        x"9",    x"8",    x"4",    x"D",    x"1",    x"A",    x"7",    x"4",
        x"D",    x"1",    x"A",    x"7",    x"4",    x"C",    x"0",    x"B",
        x"6",    x"1",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"4",    x"6",    x"8",    x"9",
        x"B",    x"D",    x"E",    x"D",    x"B",    x"9",    x"7",    x"6",
        x"4",    x"2",    x"0",    x"1",    x"2",    x"4",    x"6",    x"8",
        x"A",    x"B",    x"D",    x"E",    x"C",    x"B",    x"9",    x"7",
        x"5",    x"3",    x"2",    x"0",    x"1",    x"3",    x"4",    x"6",
        x"8",    x"A",    x"C",    x"D",    x"E",    x"C",    x"A",    x"9",
        x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",    x"5",
        x"7",    x"8",    x"A",    x"C",    x"E",    x"E",    x"C",    x"A",
        x"8",    x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",
        x"5",    x"7",    x"9",    x"A",    x"C",    x"E",    x"D",    x"C",
        x"A",    x"8",    x"6",    x"5",    x"6",    x"8",    x"C",    x"C",
        x"8",    x"4",    x"0",    x"4",    x"9",    x"D",    x"B",    x"7",
        x"2",    x"1",    x"6",    x"A",    x"E",    x"A",    x"6",    x"1",
        x"2",    x"7",    x"B",    x"D",    x"9",    x"5",    x"0",    x"3",
        x"8",    x"C",    x"C",    x"8",    x"3",    x"0",    x"5",    x"9",
        x"D",    x"B",    x"7",    x"2",    x"1",    x"6",    x"A",    x"E",
        x"A",    x"6",    x"1",    x"2",    x"7",    x"B",    x"D",    x"9",
        x"4",    x"0",    x"4",    x"8",    x"D",    x"C",    x"8",    x"3",
        x"0",    x"5",    x"9",    x"E",    x"B",    x"6",    x"0",    x"5",
        x"B",    x"C",    x"6",    x"0",    x"5",    x"B",    x"C",    x"6",
        x"0",    x"5",    x"B",    x"C",    x"6",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",
        x"A",    x"4",    x"1",    x"7",    x"D",    x"A",    x"4",    x"1",
        x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",    x"A",
        x"4",    x"2",    x"C",    x"8",    x"0",    x"9",    x"B",    x"2",
        x"6",    x"E",    x"5",    x"3",    x"C",    x"8",    x"0",    x"9",
        x"B",    x"2",    x"6",    x"F",    x"6",    x"3",    x"C",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"2",    x"B",    x"9",    x"0",    x"8",    x"C",    x"3",
        x"5",    x"E",    x"6",    x"2",    x"B",    x"9",    x"0",    x"8",
        x"C",    x"3",    x"5",    x"E",    x"6",    x"2",    x"B",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"9",    x"0",    x"C",    x"5",    x"6",    x"B",    x"0",
        x"C",    x"5",    x"6",    x"B",    x"1",    x"D",    x"4",    x"7",
        x"A",    x"1",    x"D",    x"4",    x"7",    x"A",    x"2",    x"E",
        x"3",    x"8",    x"9",    x"2",    x"E",    x"3",    x"8",    x"9",
        x"3",    x"E",    x"2",    x"9",    x"8",    x"3",    x"E",    x"2",
        x"9",    x"8",    x"4",    x"D",    x"1",    x"A",    x"7",    x"4",
        x"D",    x"1",    x"A",    x"7",    x"4",    x"C",    x"0",    x"B",
        x"6",    x"1",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"1",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"4",    x"6",    x"8",    x"9",
        x"B",    x"D",    x"E",    x"D",    x"B",    x"9",    x"7",    x"6",
        x"4",    x"2",    x"0",    x"1",    x"2",    x"4",    x"6",    x"8",
        x"A",    x"B",    x"D",    x"E",    x"C",    x"B",    x"9",    x"7",
        x"5",    x"3",    x"2",    x"0",    x"1",    x"3",    x"4",    x"6",
        x"8",    x"A",    x"C",    x"D",    x"E",    x"C",    x"A",    x"9",
        x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",    x"5",
        x"7",    x"8",    x"A",    x"C",    x"E",    x"E",    x"C",    x"A",
        x"8",    x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",
        x"5",    x"7",    x"9",    x"A",    x"C",    x"E",    x"D",    x"C",
        x"A",    x"8",    x"6",    x"5",    x"6",    x"8",    x"C",    x"C",
        x"8",    x"4",    x"0",    x"4",    x"9",    x"D",    x"B",    x"7",
        x"2",    x"1",    x"6",    x"A",    x"E",    x"A",    x"6",    x"1",
        x"2",    x"7",    x"B",    x"D",    x"9",    x"5",    x"0",    x"3",
        x"8",    x"C",    x"C",    x"8",    x"3",    x"0",    x"5",    x"9",
        x"D",    x"B",    x"7",    x"2",    x"1",    x"6",    x"A",    x"E",
        x"A",    x"6",    x"1",    x"2",    x"7",    x"B",    x"D",    x"9",
        x"4",    x"0",    x"4",    x"8",    x"D",    x"C",    x"8",    x"3",
        x"0",    x"5",    x"9",    x"E",    x"B",    x"6",    x"0",    x"5",
        x"B",    x"C",    x"6",    x"0",    x"5",    x"B",    x"C",    x"6",
        x"0",    x"5",    x"B",    x"C",    x"6",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",
        x"A",    x"4",    x"1",    x"7",    x"D",    x"A",    x"4",    x"1",
        x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",    x"A",
        x"4",    x"2",    x"C",    x"8",    x"0",    x"9",    x"B",    x"2",
        x"6",    x"E",    x"5",    x"3",    x"C",    x"8",    x"0",    x"9",
        x"B",    x"2",    x"6",    x"F",    x"6",    x"3",    x"C",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"2",    x"B",    x"9",    x"0",    x"8",    x"C",    x"3",
        x"5",    x"E",    x"6",    x"2",    x"B",    x"9",    x"0",    x"8",
        x"C",    x"3",    x"5",    x"E",    x"6",    x"2",    x"B",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"9",    x"0",    x"C",    x"5",    x"6",    x"B",    x"0",
        x"C",    x"5",    x"6",    x"B",    x"1",    x"D",    x"4",    x"7",
        x"A",    x"1",    x"D",    x"4",    x"7",    x"A",    x"2",    x"E",
        x"3",    x"8",    x"9",    x"2",    x"E",    x"3",    x"8",    x"9",
        x"3",    x"E",    x"2",    x"9",    x"8",    x"3",    x"E",    x"2",
        x"9",    x"8",    x"4",    x"D",    x"1",    x"A",    x"7",    x"4",
        x"D",    x"1",    x"A",    x"7",    x"4",    x"C",    x"0",    x"B",
        x"6",    x"1",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"1",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"4",    x"6",    x"8",    x"9",
        x"B",    x"D",    x"E",    x"D",    x"B",    x"9",    x"7",    x"6",
        x"4",    x"2",    x"0",    x"1",    x"2",    x"4",    x"6",    x"8",
        x"A",    x"B",    x"D",    x"E",    x"C",    x"B",    x"9",    x"7",
        x"5",    x"3",    x"2",    x"0",    x"1",    x"3",    x"4",    x"6",
        x"8",    x"A",    x"C",    x"D",    x"E",    x"C",    x"A",    x"9",
        x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",    x"5",
        x"7",    x"8",    x"A",    x"C",    x"E",    x"E",    x"C",    x"A",
        x"8",    x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",
        x"5",    x"7",    x"9",    x"A",    x"C",    x"E",    x"D",    x"C",
        x"A",    x"8",    x"6",    x"5",    x"6",    x"8",    x"C",    x"C",
        x"8",    x"4",    x"0",    x"4",    x"9",    x"D",    x"B",    x"7",
        x"2",    x"1",    x"6",    x"A",    x"E",    x"A",    x"6",    x"1",
        x"2",    x"7",    x"B",    x"D",    x"9",    x"5",    x"0",    x"3",
        x"8",    x"C",    x"C",    x"8",    x"3",    x"0",    x"5",    x"9",
        x"D",    x"B",    x"7",    x"2",    x"1",    x"6",    x"A",    x"E",
        x"A",    x"6",    x"1",    x"2",    x"7",    x"B",    x"D",    x"9",
        x"4",    x"0",    x"4",    x"8",    x"D",    x"C",    x"8",    x"3",
        x"0",    x"5",    x"9",    x"E",    x"B",    x"6",    x"0",    x"5",
        x"B",    x"C",    x"6",    x"0",    x"5",    x"B",    x"C",    x"6",
        x"0",    x"5",    x"B",    x"C",    x"6",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",
        x"A",    x"4",    x"1",    x"7",    x"D",    x"A",    x"4",    x"1",
        x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",    x"A",
        x"4",    x"2",    x"C",    x"8",    x"0",    x"9",    x"B",    x"2",
        x"6",    x"E",    x"5",    x"3",    x"C",    x"8",    x"0",    x"9",
        x"B",    x"2",    x"6",    x"F",    x"6",    x"3",    x"C",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"2",    x"B",    x"9",    x"0",    x"8",    x"C",    x"3",
        x"5",    x"E",    x"6",    x"2",    x"B",    x"9",    x"0",    x"8",
        x"C",    x"3",    x"5",    x"E",    x"6",    x"2",    x"B",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"9",    x"0",    x"C",    x"5",    x"6",    x"B",    x"0",
        x"C",    x"5",    x"6",    x"B",    x"1",    x"D",    x"4",    x"7",
        x"A",    x"1",    x"D",    x"4",    x"7",    x"A",    x"2",    x"E",
        x"3",    x"8",    x"9",    x"2",    x"E",    x"3",    x"8",    x"9",
        x"3",    x"E",    x"2",    x"9",    x"8",    x"3",    x"E",    x"2",
        x"9",    x"8",    x"4",    x"D",    x"1",    x"A",    x"7",    x"4",
        x"D",    x"1",    x"A",    x"7",    x"4",    x"C",    x"0",    x"B",
        x"6",    x"1",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"4",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"4",    x"6",    x"8",    x"9",
        x"B",    x"D",    x"E",    x"D",    x"B",    x"9",    x"7",    x"6",
        x"4",    x"2",    x"0",    x"1",    x"2",    x"4",    x"6",    x"8",
        x"A",    x"B",    x"D",    x"E",    x"C",    x"B",    x"9",    x"7",
        x"5",    x"3",    x"2",    x"0",    x"1",    x"3",    x"4",    x"6",
        x"8",    x"A",    x"C",    x"D",    x"E",    x"C",    x"A",    x"9",
        x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",    x"5",
        x"7",    x"8",    x"A",    x"C",    x"E",    x"E",    x"C",    x"A",
        x"8",    x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",
        x"5",    x"7",    x"9",    x"A",    x"C",    x"E",    x"D",    x"C",
        x"A",    x"8",    x"6",    x"5",    x"6",    x"8",    x"C",    x"C",
        x"8",    x"4",    x"0",    x"4",    x"9",    x"D",    x"B",    x"7",
        x"2",    x"1",    x"6",    x"A",    x"E",    x"A",    x"6",    x"1",
        x"2",    x"7",    x"B",    x"D",    x"9",    x"5",    x"0",    x"3",
        x"8",    x"C",    x"C",    x"8",    x"3",    x"0",    x"5",    x"9",
        x"D",    x"B",    x"7",    x"2",    x"1",    x"6",    x"A",    x"E",
        x"A",    x"6",    x"1",    x"2",    x"7",    x"B",    x"D",    x"9",
        x"4",    x"0",    x"4",    x"8",    x"D",    x"C",    x"8",    x"3",
        x"0",    x"5",    x"9",    x"E",    x"B",    x"6",    x"0",    x"5",
        x"B",    x"C",    x"6",    x"0",    x"5",    x"B",    x"C",    x"6",
        x"0",    x"5",    x"B",    x"C",    x"6",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",
        x"A",    x"4",    x"1",    x"7",    x"D",    x"A",    x"4",    x"1",
        x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",    x"A",
        x"4",    x"2",    x"C",    x"8",    x"0",    x"9",    x"B",    x"2",
        x"6",    x"E",    x"5",    x"3",    x"C",    x"8",    x"0",    x"9",
        x"B",    x"2",    x"6",    x"F",    x"6",    x"3",    x"C",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"2",    x"B",    x"9",    x"0",    x"8",    x"C",    x"3",
        x"5",    x"E",    x"6",    x"2",    x"B",    x"9",    x"0",    x"8",
        x"C",    x"3",    x"5",    x"E",    x"6",    x"2",    x"B",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"9",    x"0",    x"C",    x"5",    x"6",    x"B",    x"0",
        x"C",    x"5",    x"6",    x"B",    x"1",    x"D",    x"4",    x"7",
        x"A",    x"1",    x"D",    x"4",    x"7",    x"A",    x"2",    x"E",
        x"3",    x"8",    x"9",    x"2",    x"E",    x"3",    x"8",    x"9",
        x"3",    x"E",    x"2",    x"9",    x"8",    x"3",    x"E",    x"2",
        x"9",    x"8",    x"4",    x"D",    x"1",    x"A",    x"7",    x"4",
        x"D",    x"1",    x"A",    x"7",    x"4",    x"C",    x"0",    x"B",
        x"6",    x"1",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"4",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"5",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"4",    x"6",    x"8",    x"9",
        x"B",    x"D",    x"E",    x"D",    x"B",    x"9",    x"7",    x"6",
        x"4",    x"2",    x"0",    x"1",    x"2",    x"4",    x"6",    x"8",
        x"A",    x"B",    x"D",    x"E",    x"C",    x"B",    x"9",    x"7",
        x"5",    x"3",    x"2",    x"0",    x"1",    x"3",    x"4",    x"6",
        x"8",    x"A",    x"C",    x"D",    x"E",    x"C",    x"A",    x"9",
        x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",    x"5",
        x"7",    x"8",    x"A",    x"C",    x"E",    x"E",    x"C",    x"A",
        x"8",    x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",
        x"5",    x"7",    x"9",    x"A",    x"C",    x"E",    x"D",    x"C",
        x"A",    x"8",    x"6",    x"5",    x"6",    x"8",    x"C",    x"C",
        x"8",    x"4",    x"0",    x"4",    x"9",    x"D",    x"B",    x"7",
        x"2",    x"1",    x"6",    x"A",    x"E",    x"A",    x"6",    x"1",
        x"2",    x"7",    x"B",    x"D",    x"9",    x"5",    x"0",    x"3",
        x"8",    x"C",    x"C",    x"8",    x"3",    x"0",    x"5",    x"9",
        x"D",    x"B",    x"7",    x"2",    x"1",    x"6",    x"A",    x"E",
        x"A",    x"6",    x"1",    x"2",    x"7",    x"B",    x"D",    x"9",
        x"4",    x"0",    x"4",    x"8",    x"D",    x"C",    x"8",    x"3",
        x"0",    x"5",    x"9",    x"E",    x"B",    x"6",    x"0",    x"5",
        x"B",    x"C",    x"6",    x"0",    x"5",    x"B",    x"C",    x"6",
        x"0",    x"5",    x"B",    x"C",    x"6",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",
        x"A",    x"4",    x"1",    x"7",    x"D",    x"A",    x"4",    x"1",
        x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",    x"A",
        x"4",    x"2",    x"C",    x"8",    x"0",    x"9",    x"B",    x"2",
        x"6",    x"E",    x"5",    x"3",    x"C",    x"8",    x"0",    x"9",
        x"B",    x"2",    x"6",    x"F",    x"6",    x"3",    x"C",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"2",    x"B",    x"9",    x"0",    x"8",    x"C",    x"3",
        x"5",    x"E",    x"6",    x"2",    x"B",    x"9",    x"0",    x"8",
        x"C",    x"3",    x"5",    x"E",    x"6",    x"2",    x"B",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"9",    x"0",    x"C",    x"5",    x"6",    x"B",    x"0",
        x"C",    x"5",    x"6",    x"B",    x"1",    x"D",    x"4",    x"7",
        x"A",    x"1",    x"D",    x"4",    x"7",    x"A",    x"2",    x"E",
        x"3",    x"8",    x"9",    x"2",    x"E",    x"3",    x"8",    x"9",
        x"3",    x"E",    x"2",    x"9",    x"8",    x"3",    x"E",    x"2",
        x"9",    x"8",    x"4",    x"D",    x"1",    x"A",    x"7",    x"4",
        x"D",    x"1",    x"A",    x"7",    x"4",    x"C",    x"0",    x"B",
        x"6",    x"1",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"5",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"6",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"4",    x"6",    x"8",    x"9",
        x"B",    x"D",    x"E",    x"D",    x"B",    x"9",    x"7",    x"6",
        x"4",    x"2",    x"0",    x"1",    x"2",    x"4",    x"6",    x"8",
        x"A",    x"B",    x"D",    x"E",    x"C",    x"B",    x"9",    x"7",
        x"5",    x"3",    x"2",    x"0",    x"1",    x"3",    x"4",    x"6",
        x"8",    x"A",    x"C",    x"D",    x"E",    x"C",    x"A",    x"9",
        x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",    x"5",
        x"7",    x"8",    x"A",    x"C",    x"E",    x"E",    x"C",    x"A",
        x"8",    x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",
        x"5",    x"7",    x"9",    x"A",    x"C",    x"E",    x"D",    x"C",
        x"A",    x"8",    x"6",    x"5",    x"6",    x"8",    x"C",    x"C",
        x"8",    x"4",    x"0",    x"4",    x"9",    x"D",    x"B",    x"7",
        x"2",    x"1",    x"6",    x"A",    x"E",    x"A",    x"6",    x"1",
        x"2",    x"7",    x"B",    x"D",    x"9",    x"5",    x"0",    x"3",
        x"8",    x"C",    x"C",    x"8",    x"3",    x"0",    x"5",    x"9",
        x"D",    x"B",    x"7",    x"2",    x"1",    x"6",    x"A",    x"E",
        x"A",    x"6",    x"1",    x"2",    x"7",    x"B",    x"D",    x"9",
        x"4",    x"0",    x"4",    x"8",    x"D",    x"C",    x"8",    x"3",
        x"0",    x"5",    x"9",    x"E",    x"B",    x"6",    x"0",    x"5",
        x"B",    x"C",    x"6",    x"0",    x"5",    x"B",    x"C",    x"6",
        x"0",    x"5",    x"B",    x"C",    x"6",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",
        x"A",    x"4",    x"1",    x"7",    x"D",    x"A",    x"4",    x"1",
        x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",    x"A",
        x"4",    x"2",    x"C",    x"8",    x"0",    x"9",    x"B",    x"2",
        x"6",    x"E",    x"5",    x"3",    x"C",    x"8",    x"0",    x"9",
        x"B",    x"2",    x"6",    x"F",    x"6",    x"3",    x"C",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"2",    x"B",    x"9",    x"0",    x"8",    x"C",    x"3",
        x"5",    x"E",    x"6",    x"2",    x"B",    x"9",    x"0",    x"8",
        x"C",    x"3",    x"5",    x"E",    x"6",    x"2",    x"B",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"9",    x"0",    x"C",    x"5",    x"6",    x"B",    x"0",
        x"C",    x"5",    x"6",    x"B",    x"1",    x"D",    x"4",    x"7",
        x"A",    x"1",    x"D",    x"4",    x"7",    x"A",    x"2",    x"E",
        x"3",    x"8",    x"9",    x"2",    x"E",    x"3",    x"8",    x"9",
        x"3",    x"E",    x"2",    x"9",    x"8",    x"3",    x"E",    x"2",
        x"9",    x"8",    x"4",    x"D",    x"1",    x"A",    x"7",    x"4",
        x"D",    x"1",    x"A",    x"7",    x"4",    x"C",    x"0",    x"B",
        x"6",    x"1",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"4",    x"6",    x"8",    x"9",
        x"B",    x"D",    x"E",    x"D",    x"B",    x"9",    x"7",    x"6",
        x"4",    x"2",    x"0",    x"1",    x"2",    x"4",    x"6",    x"8",
        x"A",    x"B",    x"D",    x"E",    x"C",    x"B",    x"9",    x"7",
        x"5",    x"3",    x"2",    x"0",    x"1",    x"3",    x"4",    x"6",
        x"8",    x"A",    x"C",    x"D",    x"E",    x"C",    x"A",    x"9",
        x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",    x"5",
        x"7",    x"8",    x"A",    x"C",    x"E",    x"E",    x"C",    x"A",
        x"8",    x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",
        x"5",    x"7",    x"9",    x"A",    x"C",    x"E",    x"D",    x"C",
        x"A",    x"8",    x"6",    x"5",    x"6",    x"8",    x"C",    x"C",
        x"8",    x"4",    x"0",    x"4",    x"9",    x"D",    x"B",    x"7",
        x"2",    x"1",    x"6",    x"A",    x"E",    x"A",    x"6",    x"1",
        x"2",    x"7",    x"B",    x"D",    x"9",    x"5",    x"0",    x"3",
        x"8",    x"C",    x"C",    x"8",    x"3",    x"0",    x"5",    x"9",
        x"D",    x"B",    x"7",    x"2",    x"1",    x"6",    x"A",    x"E",
        x"A",    x"6",    x"1",    x"2",    x"7",    x"B",    x"D",    x"9",
        x"4",    x"0",    x"4",    x"8",    x"D",    x"C",    x"8",    x"3",
        x"0",    x"5",    x"9",    x"E",    x"B",    x"6",    x"0",    x"5",
        x"B",    x"C",    x"6",    x"0",    x"5",    x"B",    x"C",    x"6",
        x"0",    x"5",    x"B",    x"C",    x"6",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",
        x"A",    x"4",    x"1",    x"7",    x"D",    x"A",    x"4",    x"1",
        x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",    x"A",
        x"4",    x"2",    x"C",    x"8",    x"0",    x"9",    x"B",    x"2",
        x"6",    x"E",    x"5",    x"3",    x"C",    x"8",    x"0",    x"9",
        x"B",    x"2",    x"6",    x"F",    x"6",    x"3",    x"C",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"2",    x"B",    x"9",    x"0",    x"8",    x"C",    x"3",
        x"5",    x"E",    x"6",    x"2",    x"B",    x"9",    x"0",    x"8",
        x"C",    x"3",    x"5",    x"E",    x"6",    x"2",    x"B",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"9",    x"0",    x"C",    x"5",    x"6",    x"B",    x"0",
        x"C",    x"5",    x"6",    x"B",    x"1",    x"D",    x"4",    x"7",
        x"A",    x"1",    x"D",    x"4",    x"7",    x"A",    x"2",    x"E",
        x"3",    x"8",    x"9",    x"2",    x"E",    x"3",    x"8",    x"9",
        x"3",    x"E",    x"2",    x"9",    x"8",    x"3",    x"E",    x"2",
        x"9",    x"8",    x"4",    x"D",    x"1",    x"A",    x"7",    x"4",
        x"D",    x"1",    x"A",    x"7",    x"4",    x"C",    x"0",    x"B",
        x"6",    x"1",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"4",    x"6",    x"8",    x"9",
        x"B",    x"D",    x"E",    x"D",    x"B",    x"9",    x"7",    x"6",
        x"4",    x"2",    x"0",    x"1",    x"2",    x"4",    x"6",    x"8",
        x"A",    x"B",    x"D",    x"E",    x"C",    x"B",    x"9",    x"7",
        x"5",    x"3",    x"2",    x"0",    x"1",    x"3",    x"4",    x"6",
        x"8",    x"A",    x"C",    x"D",    x"E",    x"C",    x"A",    x"9",
        x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",    x"5",
        x"7",    x"8",    x"A",    x"C",    x"E",    x"E",    x"C",    x"A",
        x"8",    x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",
        x"5",    x"7",    x"9",    x"A",    x"C",    x"E",    x"D",    x"C",
        x"A",    x"8",    x"6",    x"5",    x"6",    x"8",    x"C",    x"C",
        x"8",    x"4",    x"0",    x"4",    x"9",    x"D",    x"B",    x"7",
        x"2",    x"1",    x"6",    x"A",    x"E",    x"A",    x"6",    x"1",
        x"2",    x"7",    x"B",    x"D",    x"9",    x"5",    x"0",    x"3",
        x"8",    x"C",    x"C",    x"8",    x"3",    x"0",    x"5",    x"9",
        x"D",    x"B",    x"7",    x"2",    x"1",    x"6",    x"A",    x"E",
        x"A",    x"6",    x"1",    x"2",    x"7",    x"B",    x"D",    x"9",
        x"4",    x"0",    x"4",    x"8",    x"D",    x"C",    x"8",    x"3",
        x"0",    x"5",    x"9",    x"E",    x"B",    x"6",    x"0",    x"5",
        x"B",    x"C",    x"6",    x"0",    x"5",    x"B",    x"C",    x"6",
        x"0",    x"5",    x"B",    x"C",    x"6",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",
        x"A",    x"4",    x"1",    x"7",    x"D",    x"A",    x"4",    x"1",
        x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",    x"A",
        x"4",    x"2",    x"C",    x"8",    x"0",    x"9",    x"B",    x"2",
        x"6",    x"E",    x"5",    x"3",    x"C",    x"8",    x"0",    x"9",
        x"B",    x"2",    x"6",    x"F",    x"6",    x"3",    x"C",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"2",    x"B",    x"9",    x"0",    x"8",    x"C",    x"3",
        x"5",    x"E",    x"6",    x"2",    x"B",    x"9",    x"0",    x"8",
        x"C",    x"3",    x"5",    x"E",    x"6",    x"2",    x"B",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"9",    x"0",    x"C",    x"5",    x"6",    x"B",    x"0",
        x"C",    x"5",    x"6",    x"B",    x"1",    x"D",    x"4",    x"7",
        x"A",    x"1",    x"D",    x"4",    x"7",    x"A",    x"2",    x"E",
        x"3",    x"8",    x"9",    x"2",    x"E",    x"3",    x"8",    x"9",
        x"3",    x"E",    x"2",    x"9",    x"8",    x"3",    x"E",    x"2",
        x"9",    x"8",    x"4",    x"D",    x"1",    x"A",    x"7",    x"4",
        x"D",    x"1",    x"A",    x"7",    x"4",    x"C",    x"0",    x"B",
        x"6",    x"1",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"1",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"4",    x"6",    x"8",    x"9",
        x"B",    x"D",    x"E",    x"D",    x"B",    x"9",    x"7",    x"6",
        x"4",    x"2",    x"0",    x"1",    x"2",    x"4",    x"6",    x"8",
        x"A",    x"B",    x"D",    x"E",    x"C",    x"B",    x"9",    x"7",
        x"5",    x"3",    x"2",    x"0",    x"1",    x"3",    x"4",    x"6",
        x"8",    x"A",    x"C",    x"D",    x"E",    x"C",    x"A",    x"9",
        x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",    x"5",
        x"7",    x"8",    x"A",    x"C",    x"E",    x"E",    x"C",    x"A",
        x"8",    x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",
        x"5",    x"7",    x"9",    x"A",    x"C",    x"E",    x"D",    x"C",
        x"A",    x"8",    x"6",    x"5",    x"6",    x"8",    x"C",    x"C",
        x"8",    x"4",    x"0",    x"4",    x"9",    x"D",    x"B",    x"7",
        x"2",    x"1",    x"6",    x"A",    x"E",    x"A",    x"6",    x"1",
        x"2",    x"7",    x"B",    x"D",    x"9",    x"5",    x"0",    x"3",
        x"8",    x"C",    x"C",    x"8",    x"3",    x"0",    x"5",    x"9",
        x"D",    x"B",    x"7",    x"2",    x"1",    x"6",    x"A",    x"E",
        x"A",    x"6",    x"1",    x"2",    x"7",    x"B",    x"D",    x"9",
        x"4",    x"0",    x"4",    x"8",    x"D",    x"C",    x"8",    x"3",
        x"0",    x"5",    x"9",    x"E",    x"B",    x"6",    x"0",    x"5",
        x"B",    x"C",    x"6",    x"0",    x"5",    x"B",    x"C",    x"6",
        x"0",    x"5",    x"B",    x"C",    x"6",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",
        x"A",    x"4",    x"1",    x"7",    x"D",    x"A",    x"4",    x"1",
        x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",    x"A",
        x"4",    x"2",    x"C",    x"8",    x"0",    x"9",    x"B",    x"2",
        x"6",    x"E",    x"5",    x"3",    x"C",    x"8",    x"0",    x"9",
        x"B",    x"2",    x"6",    x"F",    x"6",    x"3",    x"C",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"2",    x"B",    x"9",    x"0",    x"8",    x"C",    x"3",
        x"5",    x"E",    x"6",    x"2",    x"B",    x"9",    x"0",    x"8",
        x"C",    x"3",    x"5",    x"E",    x"6",    x"2",    x"B",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"9",    x"0",    x"C",    x"5",    x"6",    x"B",    x"0",
        x"C",    x"5",    x"6",    x"B",    x"1",    x"D",    x"4",    x"7",
        x"A",    x"1",    x"D",    x"4",    x"7",    x"A",    x"2",    x"E",
        x"3",    x"8",    x"9",    x"2",    x"E",    x"3",    x"8",    x"9",
        x"3",    x"E",    x"2",    x"9",    x"8",    x"3",    x"E",    x"2",
        x"9",    x"8",    x"4",    x"D",    x"1",    x"A",    x"7",    x"4",
        x"D",    x"1",    x"A",    x"7",    x"4",    x"C",    x"0",    x"B",
        x"6",    x"1",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"1",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"4",    x"6",    x"8",    x"9",
        x"B",    x"D",    x"E",    x"D",    x"B",    x"9",    x"7",    x"6",
        x"4",    x"2",    x"0",    x"1",    x"2",    x"4",    x"6",    x"8",
        x"A",    x"B",    x"D",    x"E",    x"C",    x"B",    x"9",    x"7",
        x"5",    x"3",    x"2",    x"0",    x"1",    x"3",    x"4",    x"6",
        x"8",    x"A",    x"C",    x"D",    x"E",    x"C",    x"A",    x"9",
        x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",    x"5",
        x"7",    x"8",    x"A",    x"C",    x"E",    x"E",    x"C",    x"A",
        x"8",    x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",
        x"5",    x"7",    x"9",    x"A",    x"C",    x"E",    x"D",    x"C",
        x"A",    x"8",    x"6",    x"5",    x"6",    x"8",    x"C",    x"C",
        x"8",    x"4",    x"0",    x"4",    x"9",    x"D",    x"B",    x"7",
        x"2",    x"1",    x"6",    x"A",    x"E",    x"A",    x"6",    x"1",
        x"2",    x"7",    x"B",    x"D",    x"9",    x"5",    x"0",    x"3",
        x"8",    x"C",    x"C",    x"8",    x"3",    x"0",    x"5",    x"9",
        x"D",    x"B",    x"7",    x"2",    x"1",    x"6",    x"A",    x"E",
        x"A",    x"6",    x"1",    x"2",    x"7",    x"B",    x"D",    x"9",
        x"4",    x"0",    x"4",    x"8",    x"D",    x"C",    x"8",    x"3",
        x"0",    x"5",    x"9",    x"E",    x"B",    x"6",    x"0",    x"5",
        x"B",    x"C",    x"6",    x"0",    x"5",    x"B",    x"C",    x"6",
        x"0",    x"5",    x"B",    x"C",    x"6",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",
        x"A",    x"4",    x"1",    x"7",    x"D",    x"A",    x"4",    x"1",
        x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",    x"A",
        x"4",    x"2",    x"C",    x"8",    x"0",    x"9",    x"B",    x"2",
        x"6",    x"E",    x"5",    x"3",    x"C",    x"8",    x"0",    x"9",
        x"B",    x"2",    x"6",    x"F",    x"6",    x"3",    x"C",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"2",    x"B",    x"9",    x"0",    x"8",    x"C",    x"3",
        x"5",    x"E",    x"6",    x"2",    x"B",    x"9",    x"0",    x"8",
        x"C",    x"3",    x"5",    x"E",    x"6",    x"2",    x"B",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"9",    x"0",    x"C",    x"5",    x"6",    x"B",    x"0",
        x"C",    x"5",    x"6",    x"B",    x"1",    x"D",    x"4",    x"7",
        x"A",    x"1",    x"D",    x"4",    x"7",    x"A",    x"2",    x"E",
        x"3",    x"8",    x"9",    x"2",    x"E",    x"3",    x"8",    x"9",
        x"3",    x"E",    x"2",    x"9",    x"8",    x"3",    x"E",    x"2",
        x"9",    x"8",    x"4",    x"D",    x"1",    x"A",    x"7",    x"4",
        x"D",    x"1",    x"A",    x"7",    x"4",    x"C",    x"0",    x"B",
        x"6",    x"1",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"5",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"4",    x"6",    x"8",    x"9",
        x"B",    x"D",    x"E",    x"D",    x"B",    x"9",    x"7",    x"6",
        x"4",    x"2",    x"0",    x"1",    x"2",    x"4",    x"6",    x"8",
        x"A",    x"B",    x"D",    x"E",    x"C",    x"B",    x"9",    x"7",
        x"5",    x"3",    x"2",    x"0",    x"1",    x"3",    x"4",    x"6",
        x"8",    x"A",    x"C",    x"D",    x"E",    x"C",    x"A",    x"9",
        x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",    x"5",
        x"7",    x"8",    x"A",    x"C",    x"E",    x"E",    x"C",    x"A",
        x"8",    x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",
        x"5",    x"7",    x"9",    x"A",    x"C",    x"E",    x"D",    x"C",
        x"A",    x"8",    x"6",    x"5",    x"6",    x"8",    x"C",    x"C",
        x"8",    x"4",    x"0",    x"4",    x"9",    x"D",    x"B",    x"7",
        x"2",    x"1",    x"6",    x"A",    x"E",    x"A",    x"6",    x"1",
        x"2",    x"7",    x"B",    x"D",    x"9",    x"5",    x"0",    x"3",
        x"8",    x"C",    x"C",    x"8",    x"3",    x"0",    x"5",    x"9",
        x"D",    x"B",    x"7",    x"2",    x"1",    x"6",    x"A",    x"E",
        x"A",    x"6",    x"1",    x"2",    x"7",    x"B",    x"D",    x"9",
        x"4",    x"0",    x"4",    x"8",    x"D",    x"C",    x"8",    x"3",
        x"0",    x"5",    x"9",    x"E",    x"B",    x"6",    x"0",    x"5",
        x"B",    x"C",    x"6",    x"0",    x"5",    x"B",    x"C",    x"6",
        x"0",    x"5",    x"B",    x"C",    x"6",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",
        x"A",    x"4",    x"1",    x"7",    x"D",    x"A",    x"4",    x"1",
        x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",    x"A",
        x"4",    x"2",    x"C",    x"8",    x"0",    x"9",    x"B",    x"2",
        x"6",    x"E",    x"5",    x"3",    x"C",    x"8",    x"0",    x"9",
        x"B",    x"2",    x"6",    x"F",    x"6",    x"3",    x"C",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"2",    x"B",    x"9",    x"0",    x"8",    x"C",    x"3",
        x"5",    x"E",    x"6",    x"2",    x"B",    x"9",    x"0",    x"8",
        x"C",    x"3",    x"5",    x"E",    x"6",    x"2",    x"B",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"9",    x"0",    x"C",    x"5",    x"6",    x"B",    x"0",
        x"C",    x"5",    x"6",    x"B",    x"1",    x"D",    x"4",    x"7",
        x"A",    x"1",    x"D",    x"4",    x"7",    x"A",    x"2",    x"E",
        x"3",    x"8",    x"9",    x"2",    x"E",    x"3",    x"8",    x"9",
        x"3",    x"E",    x"2",    x"9",    x"8",    x"3",    x"E",    x"2",
        x"9",    x"8",    x"4",    x"D",    x"1",    x"A",    x"7",    x"4",
        x"D",    x"1",    x"A",    x"7",    x"4",    x"C",    x"0",    x"B",
        x"6",    x"1",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"5",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"6",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"4",    x"6",    x"8",    x"9",
        x"B",    x"D",    x"E",    x"D",    x"B",    x"9",    x"7",    x"6",
        x"4",    x"2",    x"0",    x"1",    x"2",    x"4",    x"6",    x"8",
        x"A",    x"B",    x"D",    x"E",    x"C",    x"B",    x"9",    x"7",
        x"5",    x"3",    x"2",    x"0",    x"1",    x"3",    x"4",    x"6",
        x"8",    x"A",    x"C",    x"D",    x"E",    x"C",    x"A",    x"9",
        x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",    x"5",
        x"7",    x"8",    x"A",    x"C",    x"E",    x"E",    x"C",    x"A",
        x"8",    x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",
        x"5",    x"7",    x"9",    x"A",    x"C",    x"E",    x"D",    x"C",
        x"A",    x"8",    x"6",    x"5",    x"6",    x"8",    x"C",    x"C",
        x"8",    x"4",    x"0",    x"4",    x"9",    x"D",    x"B",    x"7",
        x"2",    x"1",    x"6",    x"A",    x"E",    x"A",    x"6",    x"1",
        x"2",    x"7",    x"B",    x"D",    x"9",    x"5",    x"0",    x"3",
        x"8",    x"C",    x"C",    x"8",    x"3",    x"0",    x"5",    x"9",
        x"D",    x"B",    x"7",    x"2",    x"1",    x"6",    x"A",    x"E",
        x"A",    x"6",    x"1",    x"2",    x"7",    x"B",    x"D",    x"9",
        x"4",    x"0",    x"4",    x"8",    x"D",    x"C",    x"8",    x"3",
        x"0",    x"5",    x"9",    x"E",    x"B",    x"6",    x"0",    x"5",
        x"B",    x"C",    x"6",    x"0",    x"5",    x"B",    x"C",    x"6",
        x"0",    x"5",    x"B",    x"C",    x"6",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",
        x"A",    x"4",    x"1",    x"7",    x"D",    x"A",    x"4",    x"1",
        x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",    x"A",
        x"4",    x"2",    x"C",    x"8",    x"0",    x"9",    x"B",    x"2",
        x"6",    x"E",    x"5",    x"3",    x"C",    x"8",    x"0",    x"9",
        x"B",    x"2",    x"6",    x"F",    x"6",    x"3",    x"C",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"2",    x"B",    x"9",    x"0",    x"8",    x"C",    x"3",
        x"5",    x"E",    x"6",    x"2",    x"B",    x"9",    x"0",    x"8",
        x"C",    x"3",    x"5",    x"E",    x"6",    x"2",    x"B",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"9",    x"0",    x"C",    x"5",    x"6",    x"B",    x"0",
        x"C",    x"5",    x"6",    x"B",    x"1",    x"D",    x"4",    x"7",
        x"A",    x"1",    x"D",    x"4",    x"7",    x"A",    x"2",    x"E",
        x"3",    x"8",    x"9",    x"2",    x"E",    x"3",    x"8",    x"9",
        x"3",    x"E",    x"2",    x"9",    x"8",    x"3",    x"E",    x"2",
        x"9",    x"8",    x"4",    x"D",    x"1",    x"A",    x"7",    x"4",
        x"D",    x"1",    x"A",    x"7",    x"4",    x"C",    x"0",    x"B",
        x"6",    x"1",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"4",    x"6",    x"8",    x"9",
        x"B",    x"D",    x"E",    x"D",    x"B",    x"9",    x"7",    x"6",
        x"4",    x"2",    x"0",    x"1",    x"2",    x"4",    x"6",    x"8",
        x"A",    x"B",    x"D",    x"E",    x"C",    x"B",    x"9",    x"7",
        x"5",    x"3",    x"2",    x"0",    x"1",    x"3",    x"4",    x"6",
        x"8",    x"A",    x"C",    x"D",    x"E",    x"C",    x"A",    x"9",
        x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",    x"5",
        x"7",    x"8",    x"A",    x"C",    x"E",    x"E",    x"C",    x"A",
        x"8",    x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",
        x"5",    x"7",    x"9",    x"A",    x"C",    x"E",    x"D",    x"C",
        x"A",    x"8",    x"6",    x"5",    x"6",    x"8",    x"C",    x"C",
        x"8",    x"4",    x"0",    x"4",    x"9",    x"D",    x"B",    x"7",
        x"2",    x"1",    x"6",    x"A",    x"E",    x"A",    x"6",    x"1",
        x"2",    x"7",    x"B",    x"D",    x"9",    x"5",    x"0",    x"3",
        x"8",    x"C",    x"C",    x"8",    x"3",    x"0",    x"5",    x"9",
        x"D",    x"B",    x"7",    x"2",    x"1",    x"6",    x"A",    x"E",
        x"A",    x"6",    x"1",    x"2",    x"7",    x"B",    x"D",    x"9",
        x"4",    x"0",    x"4",    x"8",    x"D",    x"C",    x"8",    x"3",
        x"0",    x"5",    x"9",    x"E",    x"B",    x"6",    x"0",    x"5",
        x"B",    x"C",    x"6",    x"0",    x"5",    x"B",    x"C",    x"6",
        x"0",    x"5",    x"B",    x"C",    x"6",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",
        x"A",    x"4",    x"1",    x"7",    x"D",    x"A",    x"4",    x"1",
        x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",    x"A",
        x"4",    x"2",    x"C",    x"8",    x"0",    x"9",    x"B",    x"2",
        x"6",    x"E",    x"5",    x"3",    x"C",    x"8",    x"0",    x"9",
        x"B",    x"2",    x"6",    x"F",    x"6",    x"3",    x"C",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"2",    x"B",    x"9",    x"0",    x"8",    x"C",    x"3",
        x"5",    x"E",    x"6",    x"2",    x"B",    x"9",    x"0",    x"8",
        x"C",    x"3",    x"5",    x"E",    x"6",    x"2",    x"B",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"9",    x"0",    x"C",    x"5",    x"6",    x"B",    x"0",
        x"C",    x"5",    x"6",    x"B",    x"1",    x"D",    x"4",    x"7",
        x"A",    x"1",    x"D",    x"4",    x"7",    x"A",    x"2",    x"E",
        x"3",    x"8",    x"9",    x"2",    x"E",    x"3",    x"8",    x"9",
        x"3",    x"E",    x"2",    x"9",    x"8",    x"3",    x"E",    x"2",
        x"9",    x"8",    x"4",    x"D",    x"1",    x"A",    x"7",    x"4",
        x"D",    x"1",    x"A",    x"7",    x"4",    x"C",    x"0",    x"B",
        x"6",    x"1",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"4",    x"6",    x"8",    x"9",
        x"B",    x"D",    x"E",    x"D",    x"B",    x"9",    x"7",    x"6",
        x"4",    x"2",    x"0",    x"1",    x"2",    x"4",    x"6",    x"8",
        x"A",    x"B",    x"D",    x"E",    x"C",    x"B",    x"9",    x"7",
        x"5",    x"3",    x"2",    x"0",    x"1",    x"3",    x"4",    x"6",
        x"8",    x"A",    x"C",    x"D",    x"E",    x"C",    x"A",    x"9",
        x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",    x"5",
        x"7",    x"8",    x"A",    x"C",    x"E",    x"E",    x"C",    x"A",
        x"8",    x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",
        x"5",    x"7",    x"9",    x"A",    x"C",    x"E",    x"D",    x"C",
        x"A",    x"8",    x"6",    x"5",    x"6",    x"8",    x"C",    x"C",
        x"8",    x"4",    x"0",    x"4",    x"9",    x"D",    x"B",    x"7",
        x"2",    x"1",    x"6",    x"A",    x"E",    x"A",    x"6",    x"1",
        x"2",    x"7",    x"B",    x"D",    x"9",    x"5",    x"0",    x"3",
        x"8",    x"C",    x"C",    x"8",    x"3",    x"0",    x"5",    x"9",
        x"D",    x"B",    x"7",    x"2",    x"1",    x"6",    x"A",    x"E",
        x"A",    x"6",    x"1",    x"2",    x"7",    x"B",    x"D",    x"9",
        x"4",    x"0",    x"4",    x"8",    x"D",    x"C",    x"8",    x"3",
        x"0",    x"5",    x"9",    x"E",    x"B",    x"6",    x"0",    x"5",
        x"B",    x"C",    x"6",    x"0",    x"5",    x"B",    x"C",    x"6",
        x"0",    x"5",    x"B",    x"C",    x"6",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",
        x"A",    x"4",    x"1",    x"7",    x"D",    x"A",    x"4",    x"1",
        x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",    x"A",
        x"4",    x"2",    x"C",    x"8",    x"0",    x"9",    x"B",    x"2",
        x"6",    x"E",    x"5",    x"3",    x"C",    x"8",    x"0",    x"9",
        x"B",    x"2",    x"6",    x"F",    x"6",    x"3",    x"C",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"2",    x"B",    x"9",    x"0",    x"8",    x"C",    x"3",
        x"5",    x"E",    x"6",    x"2",    x"B",    x"9",    x"0",    x"8",
        x"C",    x"3",    x"5",    x"E",    x"6",    x"2",    x"B",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"9",    x"0",    x"C",    x"5",    x"6",    x"B",    x"0",
        x"C",    x"5",    x"6",    x"B",    x"1",    x"D",    x"4",    x"7",
        x"A",    x"1",    x"D",    x"4",    x"7",    x"A",    x"2",    x"E",
        x"3",    x"8",    x"9",    x"2",    x"E",    x"3",    x"8",    x"9",
        x"3",    x"E",    x"2",    x"9",    x"8",    x"3",    x"E",    x"2",
        x"9",    x"8",    x"4",    x"D",    x"1",    x"A",    x"7",    x"4",
        x"D",    x"1",    x"A",    x"7",    x"4",    x"C",    x"0",    x"B",
        x"6",    x"1",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"2",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"4",    x"6",    x"8",    x"9",
        x"B",    x"D",    x"E",    x"D",    x"B",    x"9",    x"7",    x"6",
        x"4",    x"2",    x"0",    x"1",    x"2",    x"4",    x"6",    x"8",
        x"A",    x"B",    x"D",    x"E",    x"C",    x"B",    x"9",    x"7",
        x"5",    x"3",    x"2",    x"0",    x"1",    x"3",    x"4",    x"6",
        x"8",    x"A",    x"C",    x"D",    x"E",    x"C",    x"A",    x"9",
        x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",    x"5",
        x"7",    x"8",    x"A",    x"C",    x"E",    x"E",    x"C",    x"A",
        x"8",    x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",
        x"5",    x"7",    x"9",    x"A",    x"C",    x"E",    x"D",    x"C",
        x"A",    x"8",    x"6",    x"5",    x"6",    x"8",    x"C",    x"C",
        x"8",    x"4",    x"0",    x"4",    x"9",    x"D",    x"B",    x"7",
        x"2",    x"1",    x"6",    x"A",    x"E",    x"A",    x"6",    x"1",
        x"2",    x"7",    x"B",    x"D",    x"9",    x"5",    x"0",    x"3",
        x"8",    x"C",    x"C",    x"8",    x"3",    x"0",    x"5",    x"9",
        x"D",    x"B",    x"7",    x"2",    x"1",    x"6",    x"A",    x"E",
        x"A",    x"6",    x"1",    x"2",    x"7",    x"B",    x"D",    x"9",
        x"4",    x"0",    x"4",    x"8",    x"D",    x"C",    x"8",    x"3",
        x"0",    x"5",    x"9",    x"E",    x"B",    x"6",    x"0",    x"5",
        x"B",    x"C",    x"6",    x"0",    x"5",    x"B",    x"C",    x"6",
        x"0",    x"5",    x"B",    x"C",    x"6",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",
        x"A",    x"4",    x"1",    x"7",    x"D",    x"A",    x"4",    x"1",
        x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",    x"A",
        x"4",    x"2",    x"C",    x"8",    x"0",    x"9",    x"B",    x"2",
        x"6",    x"E",    x"5",    x"3",    x"C",    x"8",    x"0",    x"9",
        x"B",    x"2",    x"6",    x"F",    x"6",    x"3",    x"C",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"2",    x"B",    x"9",    x"0",    x"8",    x"C",    x"3",
        x"5",    x"E",    x"6",    x"2",    x"B",    x"9",    x"0",    x"8",
        x"C",    x"3",    x"5",    x"E",    x"6",    x"2",    x"B",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"9",    x"0",    x"C",    x"5",    x"6",    x"B",    x"0",
        x"C",    x"5",    x"6",    x"B",    x"1",    x"D",    x"4",    x"7",
        x"A",    x"1",    x"D",    x"4",    x"7",    x"A",    x"2",    x"E",
        x"3",    x"8",    x"9",    x"2",    x"E",    x"3",    x"8",    x"9",
        x"3",    x"E",    x"2",    x"9",    x"8",    x"3",    x"E",    x"2",
        x"9",    x"8",    x"4",    x"D",    x"1",    x"A",    x"7",    x"4",
        x"D",    x"1",    x"A",    x"7",    x"4",    x"C",    x"0",    x"B",
        x"6",    x"1",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"2",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"4",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"4",    x"6",    x"8",    x"9",
        x"B",    x"D",    x"E",    x"D",    x"B",    x"9",    x"7",    x"6",
        x"4",    x"2",    x"0",    x"1",    x"2",    x"4",    x"6",    x"8",
        x"A",    x"B",    x"D",    x"E",    x"C",    x"B",    x"9",    x"7",
        x"5",    x"3",    x"2",    x"0",    x"1",    x"3",    x"4",    x"6",
        x"8",    x"A",    x"C",    x"D",    x"E",    x"C",    x"A",    x"9",
        x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",    x"5",
        x"7",    x"8",    x"A",    x"C",    x"E",    x"E",    x"C",    x"A",
        x"8",    x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",
        x"5",    x"7",    x"9",    x"A",    x"C",    x"E",    x"D",    x"C",
        x"A",    x"8",    x"6",    x"5",    x"6",    x"8",    x"C",    x"C",
        x"8",    x"4",    x"0",    x"4",    x"9",    x"D",    x"B",    x"7",
        x"2",    x"1",    x"6",    x"A",    x"E",    x"A",    x"6",    x"1",
        x"2",    x"7",    x"B",    x"D",    x"9",    x"5",    x"0",    x"3",
        x"8",    x"C",    x"C",    x"8",    x"3",    x"0",    x"5",    x"9",
        x"D",    x"B",    x"7",    x"2",    x"1",    x"6",    x"A",    x"E",
        x"A",    x"6",    x"1",    x"2",    x"7",    x"B",    x"D",    x"9",
        x"4",    x"0",    x"4",    x"8",    x"D",    x"C",    x"8",    x"3",
        x"0",    x"5",    x"9",    x"E",    x"B",    x"6",    x"0",    x"5",
        x"B",    x"C",    x"6",    x"0",    x"5",    x"B",    x"C",    x"6",
        x"0",    x"5",    x"B",    x"C",    x"6",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",
        x"A",    x"4",    x"1",    x"7",    x"D",    x"A",    x"4",    x"1",
        x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",    x"A",
        x"4",    x"2",    x"C",    x"8",    x"0",    x"9",    x"B",    x"2",
        x"6",    x"E",    x"5",    x"3",    x"C",    x"8",    x"0",    x"9",
        x"B",    x"2",    x"6",    x"F",    x"6",    x"3",    x"C",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"2",    x"B",    x"9",    x"0",    x"8",    x"C",    x"3",
        x"5",    x"E",    x"6",    x"2",    x"B",    x"9",    x"0",    x"8",
        x"C",    x"3",    x"5",    x"E",    x"6",    x"2",    x"B",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"9",    x"0",    x"C",    x"5",    x"6",    x"B",    x"0",
        x"C",    x"5",    x"6",    x"B",    x"1",    x"D",    x"4",    x"7",
        x"A",    x"1",    x"D",    x"4",    x"7",    x"A",    x"2",    x"E",
        x"3",    x"8",    x"9",    x"2",    x"E",    x"3",    x"8",    x"9",
        x"3",    x"E",    x"2",    x"9",    x"8",    x"3",    x"E",    x"2",
        x"9",    x"8",    x"4",    x"D",    x"1",    x"A",    x"7",    x"4",
        x"D",    x"1",    x"A",    x"7",    x"4",    x"C",    x"0",    x"B",
        x"6",    x"1",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"4",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"5",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"4",    x"6",    x"8",    x"9",
        x"B",    x"D",    x"E",    x"D",    x"B",    x"9",    x"7",    x"6",
        x"4",    x"2",    x"0",    x"1",    x"2",    x"4",    x"6",    x"8",
        x"A",    x"B",    x"D",    x"E",    x"C",    x"B",    x"9",    x"7",
        x"5",    x"3",    x"2",    x"0",    x"1",    x"3",    x"4",    x"6",
        x"8",    x"A",    x"C",    x"D",    x"E",    x"C",    x"A",    x"9",
        x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",    x"5",
        x"7",    x"8",    x"A",    x"C",    x"E",    x"E",    x"C",    x"A",
        x"8",    x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",
        x"5",    x"7",    x"9",    x"A",    x"C",    x"E",    x"D",    x"C",
        x"A",    x"8",    x"6",    x"5",    x"6",    x"8",    x"C",    x"C",
        x"8",    x"4",    x"0",    x"4",    x"9",    x"D",    x"B",    x"7",
        x"2",    x"1",    x"6",    x"A",    x"E",    x"A",    x"6",    x"1",
        x"2",    x"7",    x"B",    x"D",    x"9",    x"5",    x"0",    x"3",
        x"8",    x"C",    x"C",    x"8",    x"3",    x"0",    x"5",    x"9",
        x"D",    x"B",    x"7",    x"2",    x"1",    x"6",    x"A",    x"E",
        x"A",    x"6",    x"1",    x"2",    x"7",    x"B",    x"D",    x"9",
        x"4",    x"0",    x"4",    x"8",    x"D",    x"C",    x"8",    x"3",
        x"0",    x"5",    x"9",    x"E",    x"B",    x"6",    x"0",    x"5",
        x"B",    x"C",    x"6",    x"0",    x"5",    x"B",    x"C",    x"6",
        x"0",    x"5",    x"B",    x"C",    x"6",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",
        x"A",    x"4",    x"1",    x"7",    x"D",    x"A",    x"4",    x"1",
        x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",    x"A",
        x"4",    x"2",    x"C",    x"8",    x"0",    x"9",    x"B",    x"2",
        x"6",    x"E",    x"5",    x"3",    x"C",    x"8",    x"0",    x"9",
        x"B",    x"2",    x"6",    x"F",    x"6",    x"3",    x"C",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"2",    x"B",    x"9",    x"0",    x"8",    x"C",    x"3",
        x"5",    x"E",    x"6",    x"2",    x"B",    x"9",    x"0",    x"8",
        x"C",    x"3",    x"5",    x"E",    x"6",    x"2",    x"B",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"9",    x"0",    x"C",    x"5",    x"6",    x"B",    x"0",
        x"C",    x"5",    x"6",    x"B",    x"1",    x"D",    x"4",    x"7",
        x"A",    x"1",    x"D",    x"4",    x"7",    x"A",    x"2",    x"E",
        x"3",    x"8",    x"9",    x"2",    x"E",    x"3",    x"8",    x"9",
        x"3",    x"E",    x"2",    x"9",    x"8",    x"3",    x"E",    x"2",
        x"9",    x"8",    x"4",    x"D",    x"1",    x"A",    x"7",    x"4",
        x"D",    x"1",    x"A",    x"7",    x"4",    x"C",    x"0",    x"B",
        x"6",    x"1",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"5",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"6",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"4",    x"6",    x"8",    x"9",
        x"B",    x"D",    x"E",    x"D",    x"B",    x"9",    x"7",    x"6",
        x"4",    x"2",    x"0",    x"1",    x"2",    x"4",    x"6",    x"8",
        x"A",    x"B",    x"D",    x"E",    x"C",    x"B",    x"9",    x"7",
        x"5",    x"3",    x"2",    x"0",    x"1",    x"3",    x"4",    x"6",
        x"8",    x"A",    x"C",    x"D",    x"E",    x"C",    x"A",    x"9",
        x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",    x"5",
        x"7",    x"8",    x"A",    x"C",    x"E",    x"E",    x"C",    x"A",
        x"8",    x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",
        x"5",    x"7",    x"9",    x"A",    x"C",    x"E",    x"D",    x"C",
        x"A",    x"8",    x"6",    x"5",    x"6",    x"8",    x"C",    x"C",
        x"8",    x"4",    x"0",    x"4",    x"9",    x"D",    x"B",    x"7",
        x"2",    x"1",    x"6",    x"A",    x"E",    x"A",    x"6",    x"1",
        x"2",    x"7",    x"B",    x"D",    x"9",    x"5",    x"0",    x"3",
        x"8",    x"C",    x"C",    x"8",    x"3",    x"0",    x"5",    x"9",
        x"D",    x"B",    x"7",    x"2",    x"1",    x"6",    x"A",    x"E",
        x"A",    x"6",    x"1",    x"2",    x"7",    x"B",    x"D",    x"9",
        x"4",    x"0",    x"4",    x"8",    x"D",    x"C",    x"8",    x"3",
        x"0",    x"5",    x"9",    x"E",    x"B",    x"6",    x"0",    x"5",
        x"B",    x"C",    x"6",    x"0",    x"5",    x"B",    x"C",    x"6",
        x"0",    x"5",    x"B",    x"C",    x"6",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",
        x"A",    x"4",    x"1",    x"7",    x"D",    x"A",    x"4",    x"1",
        x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",    x"A",
        x"4",    x"2",    x"C",    x"8",    x"0",    x"9",    x"B",    x"2",
        x"6",    x"E",    x"5",    x"3",    x"C",    x"8",    x"0",    x"9",
        x"B",    x"2",    x"6",    x"F",    x"6",    x"3",    x"C",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"2",    x"B",    x"9",    x"0",    x"8",    x"C",    x"3",
        x"5",    x"E",    x"6",    x"2",    x"B",    x"9",    x"0",    x"8",
        x"C",    x"3",    x"5",    x"E",    x"6",    x"2",    x"B",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"9",    x"0",    x"C",    x"5",    x"6",    x"B",    x"0",
        x"C",    x"5",    x"6",    x"B",    x"1",    x"D",    x"4",    x"7",
        x"A",    x"1",    x"D",    x"4",    x"7",    x"A",    x"2",    x"E",
        x"3",    x"8",    x"9",    x"2",    x"E",    x"3",    x"8",    x"9",
        x"3",    x"E",    x"2",    x"9",    x"8",    x"3",    x"E",    x"2",
        x"9",    x"8",    x"4",    x"D",    x"1",    x"A",    x"7",    x"4",
        x"D",    x"1",    x"A",    x"7",    x"4",    x"C",    x"0",    x"B",
        x"6",    x"1",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"6",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"4",    x"6",    x"8",    x"9",
        x"B",    x"D",    x"E",    x"D",    x"B",    x"9",    x"7",    x"6",
        x"4",    x"2",    x"0",    x"1",    x"2",    x"4",    x"6",    x"8",
        x"A",    x"B",    x"D",    x"E",    x"C",    x"B",    x"9",    x"7",
        x"5",    x"3",    x"2",    x"0",    x"1",    x"3",    x"4",    x"6",
        x"8",    x"A",    x"C",    x"D",    x"E",    x"C",    x"A",    x"9",
        x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",    x"5",
        x"7",    x"8",    x"A",    x"C",    x"E",    x"E",    x"C",    x"A",
        x"8",    x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",
        x"5",    x"7",    x"9",    x"A",    x"C",    x"E",    x"D",    x"C",
        x"A",    x"8",    x"6",    x"5",    x"6",    x"8",    x"C",    x"C",
        x"8",    x"4",    x"0",    x"4",    x"9",    x"D",    x"B",    x"7",
        x"2",    x"1",    x"6",    x"A",    x"E",    x"A",    x"6",    x"1",
        x"2",    x"7",    x"B",    x"D",    x"9",    x"5",    x"0",    x"3",
        x"8",    x"C",    x"C",    x"8",    x"3",    x"0",    x"5",    x"9",
        x"D",    x"B",    x"7",    x"2",    x"1",    x"6",    x"A",    x"E",
        x"A",    x"6",    x"1",    x"2",    x"7",    x"B",    x"D",    x"9",
        x"4",    x"0",    x"4",    x"8",    x"D",    x"C",    x"8",    x"3",
        x"0",    x"5",    x"9",    x"E",    x"B",    x"6",    x"0",    x"5",
        x"B",    x"C",    x"6",    x"0",    x"5",    x"B",    x"C",    x"6",
        x"0",    x"5",    x"B",    x"C",    x"6",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",
        x"A",    x"4",    x"1",    x"7",    x"D",    x"A",    x"4",    x"1",
        x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",    x"A",
        x"4",    x"2",    x"C",    x"8",    x"0",    x"9",    x"B",    x"2",
        x"6",    x"E",    x"5",    x"3",    x"C",    x"8",    x"0",    x"9",
        x"B",    x"2",    x"6",    x"F",    x"6",    x"3",    x"C",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"2",    x"B",    x"9",    x"0",    x"8",    x"C",    x"3",
        x"5",    x"E",    x"6",    x"2",    x"B",    x"9",    x"0",    x"8",
        x"C",    x"3",    x"5",    x"E",    x"6",    x"2",    x"B",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"9",    x"0",    x"C",    x"5",    x"6",    x"B",    x"0",
        x"C",    x"5",    x"6",    x"B",    x"1",    x"D",    x"4",    x"7",
        x"A",    x"1",    x"D",    x"4",    x"7",    x"A",    x"2",    x"E",
        x"3",    x"8",    x"9",    x"2",    x"E",    x"3",    x"8",    x"9",
        x"3",    x"E",    x"2",    x"9",    x"8",    x"3",    x"E",    x"2",
        x"9",    x"8",    x"4",    x"D",    x"1",    x"A",    x"7",    x"4",
        x"D",    x"1",    x"A",    x"7",    x"4",    x"C",    x"0",    x"B",
        x"6",    x"1",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"2",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"4",    x"6",    x"8",    x"9",
        x"B",    x"D",    x"E",    x"D",    x"B",    x"9",    x"7",    x"6",
        x"4",    x"2",    x"0",    x"1",    x"2",    x"4",    x"6",    x"8",
        x"A",    x"B",    x"D",    x"E",    x"C",    x"B",    x"9",    x"7",
        x"5",    x"3",    x"2",    x"0",    x"1",    x"3",    x"4",    x"6",
        x"8",    x"A",    x"C",    x"D",    x"E",    x"C",    x"A",    x"9",
        x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",    x"5",
        x"7",    x"8",    x"A",    x"C",    x"E",    x"E",    x"C",    x"A",
        x"8",    x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",
        x"5",    x"7",    x"9",    x"A",    x"C",    x"E",    x"D",    x"C",
        x"A",    x"8",    x"6",    x"5",    x"6",    x"8",    x"C",    x"C",
        x"8",    x"4",    x"0",    x"4",    x"9",    x"D",    x"B",    x"7",
        x"2",    x"1",    x"6",    x"A",    x"E",    x"A",    x"6",    x"1",
        x"2",    x"7",    x"B",    x"D",    x"9",    x"5",    x"0",    x"3",
        x"8",    x"C",    x"C",    x"8",    x"3",    x"0",    x"5",    x"9",
        x"D",    x"B",    x"7",    x"2",    x"1",    x"6",    x"A",    x"E",
        x"A",    x"6",    x"1",    x"2",    x"7",    x"B",    x"D",    x"9",
        x"4",    x"0",    x"4",    x"8",    x"D",    x"C",    x"8",    x"3",
        x"0",    x"5",    x"9",    x"E",    x"B",    x"6",    x"0",    x"5",
        x"B",    x"C",    x"6",    x"0",    x"5",    x"B",    x"C",    x"6",
        x"0",    x"5",    x"B",    x"C",    x"6",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",
        x"A",    x"4",    x"1",    x"7",    x"D",    x"A",    x"4",    x"1",
        x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",    x"A",
        x"4",    x"2",    x"C",    x"8",    x"0",    x"9",    x"B",    x"2",
        x"6",    x"E",    x"5",    x"3",    x"C",    x"8",    x"0",    x"9",
        x"B",    x"2",    x"6",    x"F",    x"6",    x"3",    x"C",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"2",    x"B",    x"9",    x"0",    x"8",    x"C",    x"3",
        x"5",    x"E",    x"6",    x"2",    x"B",    x"9",    x"0",    x"8",
        x"C",    x"3",    x"5",    x"E",    x"6",    x"2",    x"B",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"9",    x"0",    x"C",    x"5",    x"6",    x"B",    x"0",
        x"C",    x"5",    x"6",    x"B",    x"1",    x"D",    x"4",    x"7",
        x"A",    x"1",    x"D",    x"4",    x"7",    x"A",    x"2",    x"E",
        x"3",    x"8",    x"9",    x"2",    x"E",    x"3",    x"8",    x"9",
        x"3",    x"E",    x"2",    x"9",    x"8",    x"3",    x"E",    x"2",
        x"9",    x"8",    x"4",    x"D",    x"1",    x"A",    x"7",    x"4",
        x"D",    x"1",    x"A",    x"7",    x"4",    x"C",    x"0",    x"B",
        x"6",    x"1",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"4",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"4",    x"6",    x"8",    x"9",
        x"B",    x"D",    x"E",    x"D",    x"B",    x"9",    x"7",    x"6",
        x"4",    x"2",    x"0",    x"1",    x"2",    x"4",    x"6",    x"8",
        x"A",    x"B",    x"D",    x"E",    x"C",    x"B",    x"9",    x"7",
        x"5",    x"3",    x"2",    x"0",    x"1",    x"3",    x"4",    x"6",
        x"8",    x"A",    x"C",    x"D",    x"E",    x"C",    x"A",    x"9",
        x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",    x"5",
        x"7",    x"8",    x"A",    x"C",    x"E",    x"E",    x"C",    x"A",
        x"8",    x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",
        x"5",    x"7",    x"9",    x"A",    x"C",    x"E",    x"D",    x"C",
        x"A",    x"8",    x"6",    x"5",    x"6",    x"8",    x"C",    x"C",
        x"8",    x"4",    x"0",    x"4",    x"9",    x"D",    x"B",    x"7",
        x"2",    x"1",    x"6",    x"A",    x"E",    x"A",    x"6",    x"1",
        x"2",    x"7",    x"B",    x"D",    x"9",    x"5",    x"0",    x"3",
        x"8",    x"C",    x"C",    x"8",    x"3",    x"0",    x"5",    x"9",
        x"D",    x"B",    x"7",    x"2",    x"1",    x"6",    x"A",    x"E",
        x"A",    x"6",    x"1",    x"2",    x"7",    x"B",    x"D",    x"9",
        x"4",    x"0",    x"4",    x"8",    x"D",    x"C",    x"8",    x"3",
        x"0",    x"5",    x"9",    x"E",    x"B",    x"6",    x"0",    x"5",
        x"B",    x"C",    x"6",    x"0",    x"5",    x"B",    x"C",    x"6",
        x"0",    x"5",    x"B",    x"C",    x"6",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",
        x"A",    x"4",    x"1",    x"7",    x"D",    x"A",    x"4",    x"1",
        x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",    x"A",
        x"4",    x"2",    x"C",    x"8",    x"0",    x"9",    x"B",    x"2",
        x"6",    x"E",    x"5",    x"3",    x"C",    x"8",    x"0",    x"9",
        x"B",    x"2",    x"6",    x"F",    x"6",    x"3",    x"C",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"2",    x"B",    x"9",    x"0",    x"8",    x"C",    x"3",
        x"5",    x"E",    x"6",    x"2",    x"B",    x"9",    x"0",    x"8",
        x"C",    x"3",    x"5",    x"E",    x"6",    x"2",    x"B",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"9",    x"0",    x"C",    x"5",    x"6",    x"B",    x"0",
        x"C",    x"5",    x"6",    x"B",    x"1",    x"D",    x"4",    x"7",
        x"A",    x"1",    x"D",    x"4",    x"7",    x"A",    x"2",    x"E",
        x"3",    x"8",    x"9",    x"2",    x"E",    x"3",    x"8",    x"9",
        x"3",    x"E",    x"2",    x"9",    x"8",    x"3",    x"E",    x"2",
        x"9",    x"8",    x"4",    x"D",    x"1",    x"A",    x"7",    x"4",
        x"D",    x"1",    x"A",    x"7",    x"4",    x"C",    x"0",    x"B",
        x"6",    x"1",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"4",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"6",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"4",    x"6",    x"8",    x"9",
        x"B",    x"D",    x"E",    x"D",    x"B",    x"9",    x"7",    x"6",
        x"4",    x"2",    x"0",    x"1",    x"2",    x"4",    x"6",    x"8",
        x"A",    x"B",    x"D",    x"E",    x"C",    x"B",    x"9",    x"7",
        x"5",    x"3",    x"2",    x"0",    x"1",    x"3",    x"4",    x"6",
        x"8",    x"A",    x"C",    x"D",    x"E",    x"C",    x"A",    x"9",
        x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",    x"5",
        x"7",    x"8",    x"A",    x"C",    x"E",    x"E",    x"C",    x"A",
        x"8",    x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",
        x"5",    x"7",    x"9",    x"A",    x"C",    x"E",    x"D",    x"C",
        x"A",    x"8",    x"6",    x"5",    x"6",    x"8",    x"C",    x"C",
        x"8",    x"4",    x"0",    x"4",    x"9",    x"D",    x"B",    x"7",
        x"2",    x"1",    x"6",    x"A",    x"E",    x"A",    x"6",    x"1",
        x"2",    x"7",    x"B",    x"D",    x"9",    x"5",    x"0",    x"3",
        x"8",    x"C",    x"C",    x"8",    x"3",    x"0",    x"5",    x"9",
        x"D",    x"B",    x"7",    x"2",    x"1",    x"6",    x"A",    x"E",
        x"A",    x"6",    x"1",    x"2",    x"7",    x"B",    x"D",    x"9",
        x"4",    x"0",    x"4",    x"8",    x"D",    x"C",    x"8",    x"3",
        x"0",    x"5",    x"9",    x"E",    x"B",    x"6",    x"0",    x"5",
        x"B",    x"C",    x"6",    x"0",    x"5",    x"B",    x"C",    x"6",
        x"0",    x"5",    x"B",    x"C",    x"6",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",
        x"A",    x"4",    x"1",    x"7",    x"D",    x"A",    x"4",    x"1",
        x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",    x"A",
        x"4",    x"2",    x"C",    x"8",    x"0",    x"9",    x"B",    x"2",
        x"6",    x"E",    x"5",    x"3",    x"C",    x"8",    x"0",    x"9",
        x"B",    x"2",    x"6",    x"F",    x"6",    x"3",    x"C",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"2",    x"B",    x"9",    x"0",    x"8",    x"C",    x"3",
        x"5",    x"E",    x"6",    x"2",    x"B",    x"9",    x"0",    x"8",
        x"C",    x"3",    x"5",    x"E",    x"6",    x"2",    x"B",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"9",    x"0",    x"C",    x"5",    x"6",    x"B",    x"0",
        x"C",    x"5",    x"6",    x"B",    x"1",    x"D",    x"4",    x"7",
        x"A",    x"1",    x"D",    x"4",    x"7",    x"A",    x"2",    x"E",
        x"3",    x"8",    x"9",    x"2",    x"E",    x"3",    x"8",    x"9",
        x"3",    x"E",    x"2",    x"9",    x"8",    x"3",    x"E",    x"2",
        x"9",    x"8",    x"4",    x"D",    x"1",    x"A",    x"7",    x"4",
        x"D",    x"1",    x"A",    x"7",    x"4",    x"C",    x"0",    x"B",
        x"6",    x"1",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"6",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"4",    x"6",    x"8",    x"9",
        x"B",    x"D",    x"E",    x"D",    x"B",    x"9",    x"7",    x"6",
        x"4",    x"2",    x"0",    x"1",    x"2",    x"4",    x"6",    x"8",
        x"A",    x"B",    x"D",    x"E",    x"C",    x"B",    x"9",    x"7",
        x"5",    x"3",    x"2",    x"0",    x"1",    x"3",    x"4",    x"6",
        x"8",    x"A",    x"C",    x"D",    x"E",    x"C",    x"A",    x"9",
        x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",    x"5",
        x"7",    x"8",    x"A",    x"C",    x"E",    x"E",    x"C",    x"A",
        x"8",    x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",
        x"5",    x"7",    x"9",    x"A",    x"C",    x"E",    x"D",    x"C",
        x"A",    x"8",    x"6",    x"5",    x"6",    x"8",    x"C",    x"C",
        x"8",    x"4",    x"0",    x"4",    x"9",    x"D",    x"B",    x"7",
        x"2",    x"1",    x"6",    x"A",    x"E",    x"A",    x"6",    x"1",
        x"2",    x"7",    x"B",    x"D",    x"9",    x"5",    x"0",    x"3",
        x"8",    x"C",    x"C",    x"8",    x"3",    x"0",    x"5",    x"9",
        x"D",    x"B",    x"7",    x"2",    x"1",    x"6",    x"A",    x"E",
        x"A",    x"6",    x"1",    x"2",    x"7",    x"B",    x"D",    x"9",
        x"4",    x"0",    x"4",    x"8",    x"D",    x"C",    x"8",    x"3",
        x"0",    x"5",    x"9",    x"E",    x"B",    x"6",    x"0",    x"5",
        x"B",    x"C",    x"6",    x"0",    x"5",    x"B",    x"C",    x"6",
        x"0",    x"5",    x"B",    x"C",    x"6",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",
        x"A",    x"4",    x"1",    x"7",    x"D",    x"A",    x"4",    x"1",
        x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",    x"A",
        x"4",    x"2",    x"C",    x"8",    x"0",    x"9",    x"B",    x"2",
        x"6",    x"E",    x"5",    x"3",    x"C",    x"8",    x"0",    x"9",
        x"B",    x"2",    x"6",    x"F",    x"6",    x"3",    x"C",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"2",    x"B",    x"9",    x"0",    x"8",    x"C",    x"3",
        x"5",    x"E",    x"6",    x"2",    x"B",    x"9",    x"0",    x"8",
        x"C",    x"3",    x"5",    x"E",    x"6",    x"2",    x"B",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"9",    x"0",    x"C",    x"5",    x"6",    x"B",    x"0",
        x"C",    x"5",    x"6",    x"B",    x"1",    x"D",    x"4",    x"7",
        x"A",    x"1",    x"D",    x"4",    x"7",    x"A",    x"2",    x"E",
        x"3",    x"8",    x"9",    x"2",    x"E",    x"3",    x"8",    x"9",
        x"3",    x"E",    x"2",    x"9",    x"8",    x"3",    x"E",    x"2",
        x"9",    x"8",    x"4",    x"D",    x"1",    x"A",    x"7",    x"4",
        x"D",    x"1",    x"A",    x"7",    x"4",    x"C",    x"0",    x"B",
        x"6",    x"1",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"1",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"4",    x"6",    x"8",    x"9",
        x"B",    x"D",    x"E",    x"D",    x"B",    x"9",    x"7",    x"6",
        x"4",    x"2",    x"0",    x"1",    x"2",    x"4",    x"6",    x"8",
        x"A",    x"B",    x"D",    x"E",    x"C",    x"B",    x"9",    x"7",
        x"5",    x"3",    x"2",    x"0",    x"1",    x"3",    x"4",    x"6",
        x"8",    x"A",    x"C",    x"D",    x"E",    x"C",    x"A",    x"9",
        x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",    x"5",
        x"7",    x"8",    x"A",    x"C",    x"E",    x"E",    x"C",    x"A",
        x"8",    x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",
        x"5",    x"7",    x"9",    x"A",    x"C",    x"E",    x"D",    x"C",
        x"A",    x"8",    x"6",    x"5",    x"6",    x"8",    x"C",    x"C",
        x"8",    x"4",    x"0",    x"4",    x"9",    x"D",    x"B",    x"7",
        x"2",    x"1",    x"6",    x"A",    x"E",    x"A",    x"6",    x"1",
        x"2",    x"7",    x"B",    x"D",    x"9",    x"5",    x"0",    x"3",
        x"8",    x"C",    x"C",    x"8",    x"3",    x"0",    x"5",    x"9",
        x"D",    x"B",    x"7",    x"2",    x"1",    x"6",    x"A",    x"E",
        x"A",    x"6",    x"1",    x"2",    x"7",    x"B",    x"D",    x"9",
        x"4",    x"0",    x"4",    x"8",    x"D",    x"C",    x"8",    x"3",
        x"0",    x"5",    x"9",    x"E",    x"B",    x"6",    x"0",    x"5",
        x"B",    x"C",    x"6",    x"0",    x"5",    x"B",    x"C",    x"6",
        x"0",    x"5",    x"B",    x"C",    x"6",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",
        x"A",    x"4",    x"1",    x"7",    x"D",    x"A",    x"4",    x"1",
        x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",    x"A",
        x"4",    x"2",    x"C",    x"8",    x"0",    x"9",    x"B",    x"2",
        x"6",    x"E",    x"5",    x"3",    x"C",    x"8",    x"0",    x"9",
        x"B",    x"2",    x"6",    x"F",    x"6",    x"3",    x"C",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"2",    x"B",    x"9",    x"0",    x"8",    x"C",    x"3",
        x"5",    x"E",    x"6",    x"2",    x"B",    x"9",    x"0",    x"8",
        x"C",    x"3",    x"5",    x"E",    x"6",    x"2",    x"B",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"9",    x"0",    x"C",    x"5",    x"6",    x"B",    x"0",
        x"C",    x"5",    x"6",    x"B",    x"1",    x"D",    x"4",    x"7",
        x"A",    x"1",    x"D",    x"4",    x"7",    x"A",    x"2",    x"E",
        x"3",    x"8",    x"9",    x"2",    x"E",    x"3",    x"8",    x"9",
        x"3",    x"E",    x"2",    x"9",    x"8",    x"3",    x"E",    x"2",
        x"9",    x"8",    x"4",    x"D",    x"1",    x"A",    x"7",    x"4",
        x"D",    x"1",    x"A",    x"7",    x"4",    x"C",    x"0",    x"B",
        x"6",    x"1",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"1",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"3",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"4",    x"6",    x"8",    x"9",
        x"B",    x"D",    x"E",    x"D",    x"B",    x"9",    x"7",    x"6",
        x"4",    x"2",    x"0",    x"1",    x"2",    x"4",    x"6",    x"8",
        x"A",    x"B",    x"D",    x"E",    x"C",    x"B",    x"9",    x"7",
        x"5",    x"3",    x"2",    x"0",    x"1",    x"3",    x"4",    x"6",
        x"8",    x"A",    x"C",    x"D",    x"E",    x"C",    x"A",    x"9",
        x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",    x"5",
        x"7",    x"8",    x"A",    x"C",    x"E",    x"E",    x"C",    x"A",
        x"8",    x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",
        x"5",    x"7",    x"9",    x"A",    x"C",    x"E",    x"D",    x"C",
        x"A",    x"8",    x"6",    x"5",    x"6",    x"8",    x"C",    x"C",
        x"8",    x"4",    x"0",    x"4",    x"9",    x"D",    x"B",    x"7",
        x"2",    x"1",    x"6",    x"A",    x"E",    x"A",    x"6",    x"1",
        x"2",    x"7",    x"B",    x"D",    x"9",    x"5",    x"0",    x"3",
        x"8",    x"C",    x"C",    x"8",    x"3",    x"0",    x"5",    x"9",
        x"D",    x"B",    x"7",    x"2",    x"1",    x"6",    x"A",    x"E",
        x"A",    x"6",    x"1",    x"2",    x"7",    x"B",    x"D",    x"9",
        x"4",    x"0",    x"4",    x"8",    x"D",    x"C",    x"8",    x"3",
        x"0",    x"5",    x"9",    x"E",    x"B",    x"6",    x"0",    x"5",
        x"B",    x"C",    x"6",    x"0",    x"5",    x"B",    x"C",    x"6",
        x"0",    x"5",    x"B",    x"C",    x"6",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",
        x"A",    x"4",    x"1",    x"7",    x"D",    x"A",    x"4",    x"1",
        x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",    x"A",
        x"4",    x"2",    x"C",    x"8",    x"0",    x"9",    x"B",    x"2",
        x"6",    x"E",    x"5",    x"3",    x"C",    x"8",    x"0",    x"9",
        x"B",    x"2",    x"6",    x"F",    x"6",    x"3",    x"C",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"2",    x"B",    x"9",    x"0",    x"8",    x"C",    x"3",
        x"5",    x"E",    x"6",    x"2",    x"B",    x"9",    x"0",    x"8",
        x"C",    x"3",    x"5",    x"E",    x"6",    x"2",    x"B",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"9",    x"0",    x"C",    x"5",    x"6",    x"B",    x"0",
        x"C",    x"5",    x"6",    x"B",    x"1",    x"D",    x"4",    x"7",
        x"A",    x"1",    x"D",    x"4",    x"7",    x"A",    x"2",    x"E",
        x"3",    x"8",    x"9",    x"2",    x"E",    x"3",    x"8",    x"9",
        x"3",    x"E",    x"2",    x"9",    x"8",    x"3",    x"E",    x"2",
        x"9",    x"8",    x"4",    x"D",    x"1",    x"A",    x"7",    x"4",
        x"D",    x"1",    x"A",    x"7",    x"4",    x"C",    x"0",    x"B",
        x"6",    x"1",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"4",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"5",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"4",    x"6",    x"8",    x"9",
        x"B",    x"D",    x"E",    x"D",    x"B",    x"9",    x"7",    x"6",
        x"4",    x"2",    x"0",    x"1",    x"2",    x"4",    x"6",    x"8",
        x"A",    x"B",    x"D",    x"E",    x"C",    x"B",    x"9",    x"7",
        x"5",    x"3",    x"2",    x"0",    x"1",    x"3",    x"4",    x"6",
        x"8",    x"A",    x"C",    x"D",    x"E",    x"C",    x"A",    x"9",
        x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",    x"5",
        x"7",    x"8",    x"A",    x"C",    x"E",    x"E",    x"C",    x"A",
        x"8",    x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",
        x"5",    x"7",    x"9",    x"A",    x"C",    x"E",    x"D",    x"C",
        x"A",    x"8",    x"6",    x"5",    x"6",    x"8",    x"C",    x"C",
        x"8",    x"4",    x"0",    x"4",    x"9",    x"D",    x"B",    x"7",
        x"2",    x"1",    x"6",    x"A",    x"E",    x"A",    x"6",    x"1",
        x"2",    x"7",    x"B",    x"D",    x"9",    x"5",    x"0",    x"3",
        x"8",    x"C",    x"C",    x"8",    x"3",    x"0",    x"5",    x"9",
        x"D",    x"B",    x"7",    x"2",    x"1",    x"6",    x"A",    x"E",
        x"A",    x"6",    x"1",    x"2",    x"7",    x"B",    x"D",    x"9",
        x"4",    x"0",    x"4",    x"8",    x"D",    x"C",    x"8",    x"3",
        x"0",    x"5",    x"9",    x"E",    x"B",    x"6",    x"0",    x"5",
        x"B",    x"C",    x"6",    x"0",    x"5",    x"B",    x"C",    x"6",
        x"0",    x"5",    x"B",    x"C",    x"6",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",
        x"A",    x"4",    x"1",    x"7",    x"D",    x"A",    x"4",    x"1",
        x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",    x"A",
        x"4",    x"2",    x"C",    x"8",    x"0",    x"9",    x"B",    x"2",
        x"6",    x"E",    x"5",    x"3",    x"C",    x"8",    x"0",    x"9",
        x"B",    x"2",    x"6",    x"F",    x"6",    x"3",    x"C",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"2",    x"B",    x"9",    x"0",    x"8",    x"C",    x"3",
        x"5",    x"E",    x"6",    x"2",    x"B",    x"9",    x"0",    x"8",
        x"C",    x"3",    x"5",    x"E",    x"6",    x"2",    x"B",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"9",    x"0",    x"C",    x"5",    x"6",    x"B",    x"0",
        x"C",    x"5",    x"6",    x"B",    x"1",    x"D",    x"4",    x"7",
        x"A",    x"1",    x"D",    x"4",    x"7",    x"A",    x"2",    x"E",
        x"3",    x"8",    x"9",    x"2",    x"E",    x"3",    x"8",    x"9",
        x"3",    x"E",    x"2",    x"9",    x"8",    x"3",    x"E",    x"2",
        x"9",    x"8",    x"4",    x"D",    x"1",    x"A",    x"7",    x"4",
        x"D",    x"1",    x"A",    x"7",    x"4",    x"C",    x"0",    x"B",
        x"6",    x"1",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"6",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"D",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"C",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"9",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"4",    x"6",    x"8",    x"9",
        x"B",    x"D",    x"E",    x"D",    x"B",    x"9",    x"7",    x"6",
        x"4",    x"2",    x"0",    x"1",    x"2",    x"4",    x"6",    x"8",
        x"A",    x"B",    x"D",    x"E",    x"C",    x"B",    x"9",    x"7",
        x"5",    x"3",    x"2",    x"0",    x"1",    x"3",    x"4",    x"6",
        x"8",    x"A",    x"C",    x"D",    x"E",    x"C",    x"A",    x"9",
        x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",    x"5",
        x"7",    x"8",    x"A",    x"C",    x"E",    x"E",    x"C",    x"A",
        x"8",    x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",
        x"5",    x"7",    x"9",    x"A",    x"C",    x"E",    x"D",    x"C",
        x"A",    x"8",    x"6",    x"5",    x"6",    x"8",    x"C",    x"C",
        x"8",    x"4",    x"0",    x"4",    x"9",    x"D",    x"B",    x"7",
        x"2",    x"1",    x"6",    x"A",    x"E",    x"A",    x"6",    x"1",
        x"2",    x"7",    x"B",    x"D",    x"9",    x"5",    x"0",    x"3",
        x"8",    x"C",    x"C",    x"8",    x"3",    x"0",    x"5",    x"9",
        x"D",    x"B",    x"7",    x"2",    x"1",    x"6",    x"A",    x"E",
        x"A",    x"6",    x"1",    x"2",    x"7",    x"B",    x"D",    x"9",
        x"4",    x"0",    x"4",    x"8",    x"D",    x"C",    x"8",    x"3",
        x"0",    x"5",    x"9",    x"E",    x"B",    x"6",    x"0",    x"5",
        x"B",    x"C",    x"6",    x"0",    x"5",    x"B",    x"C",    x"6",
        x"0",    x"5",    x"B",    x"C",    x"6",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",
        x"A",    x"4",    x"1",    x"7",    x"D",    x"A",    x"4",    x"1",
        x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",    x"A",
        x"4",    x"2",    x"C",    x"8",    x"0",    x"9",    x"B",    x"2",
        x"6",    x"E",    x"5",    x"3",    x"C",    x"8",    x"0",    x"9",
        x"B",    x"2",    x"6",    x"F",    x"6",    x"3",    x"C",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"2",    x"B",    x"9",    x"0",    x"8",    x"C",    x"3",
        x"5",    x"E",    x"6",    x"2",    x"B",    x"9",    x"0",    x"8",
        x"C",    x"3",    x"5",    x"E",    x"6",    x"2",    x"B",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"9",    x"0",    x"C",    x"5",    x"6",    x"B",    x"0",
        x"C",    x"5",    x"6",    x"B",    x"1",    x"D",    x"4",    x"7",
        x"A",    x"1",    x"D",    x"4",    x"7",    x"A",    x"2",    x"E",
        x"3",    x"8",    x"9",    x"2",    x"E",    x"3",    x"8",    x"9",
        x"3",    x"E",    x"2",    x"9",    x"8",    x"3",    x"E",    x"2",
        x"9",    x"8",    x"4",    x"D",    x"1",    x"A",    x"7",    x"4",
        x"D",    x"1",    x"A",    x"7",    x"4",    x"C",    x"0",    x"B",
        x"6",    x"1",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"9",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"C",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"D",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"E",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"4",    x"6",    x"8",    x"9",
        x"B",    x"D",    x"E",    x"D",    x"B",    x"9",    x"7",    x"6",
        x"4",    x"2",    x"0",    x"1",    x"2",    x"4",    x"6",    x"8",
        x"A",    x"B",    x"D",    x"E",    x"C",    x"B",    x"9",    x"7",
        x"5",    x"3",    x"2",    x"0",    x"1",    x"3",    x"4",    x"6",
        x"8",    x"A",    x"C",    x"D",    x"E",    x"C",    x"A",    x"9",
        x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",    x"5",
        x"7",    x"8",    x"A",    x"C",    x"E",    x"E",    x"C",    x"A",
        x"8",    x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",
        x"5",    x"7",    x"9",    x"A",    x"C",    x"E",    x"D",    x"C",
        x"A",    x"8",    x"6",    x"5",    x"6",    x"8",    x"C",    x"C",
        x"8",    x"4",    x"0",    x"4",    x"9",    x"D",    x"B",    x"7",
        x"2",    x"1",    x"6",    x"A",    x"E",    x"A",    x"6",    x"1",
        x"2",    x"7",    x"B",    x"D",    x"9",    x"5",    x"0",    x"3",
        x"8",    x"C",    x"C",    x"8",    x"3",    x"0",    x"5",    x"9",
        x"D",    x"B",    x"7",    x"2",    x"1",    x"6",    x"A",    x"E",
        x"A",    x"6",    x"1",    x"2",    x"7",    x"B",    x"D",    x"9",
        x"4",    x"0",    x"4",    x"8",    x"D",    x"C",    x"8",    x"3",
        x"0",    x"5",    x"9",    x"E",    x"B",    x"6",    x"0",    x"5",
        x"B",    x"C",    x"6",    x"0",    x"5",    x"B",    x"C",    x"6",
        x"0",    x"5",    x"B",    x"C",    x"6",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",
        x"A",    x"4",    x"1",    x"7",    x"D",    x"A",    x"4",    x"1",
        x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",    x"A",
        x"4",    x"2",    x"C",    x"8",    x"0",    x"9",    x"B",    x"2",
        x"6",    x"E",    x"5",    x"3",    x"C",    x"8",    x"0",    x"9",
        x"B",    x"2",    x"6",    x"F",    x"6",    x"3",    x"C",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"2",    x"B",    x"9",    x"0",    x"8",    x"C",    x"3",
        x"5",    x"E",    x"6",    x"2",    x"B",    x"9",    x"0",    x"8",
        x"C",    x"3",    x"5",    x"E",    x"6",    x"2",    x"B",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"9",    x"0",    x"C",    x"5",    x"6",    x"B",    x"0",
        x"C",    x"5",    x"6",    x"B",    x"1",    x"D",    x"4",    x"7",
        x"A",    x"1",    x"D",    x"4",    x"7",    x"A",    x"2",    x"E",
        x"3",    x"8",    x"9",    x"2",    x"E",    x"3",    x"8",    x"9",
        x"3",    x"E",    x"2",    x"9",    x"8",    x"3",    x"E",    x"2",
        x"9",    x"8",    x"4",    x"D",    x"1",    x"A",    x"7",    x"4",
        x"D",    x"1",    x"A",    x"7",    x"4",    x"C",    x"0",    x"B",
        x"6",    x"1",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"E",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"3",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"4",    x"6",    x"8",    x"9",
        x"B",    x"D",    x"E",    x"D",    x"B",    x"9",    x"7",    x"6",
        x"4",    x"2",    x"0",    x"1",    x"2",    x"4",    x"6",    x"8",
        x"A",    x"B",    x"D",    x"E",    x"C",    x"B",    x"9",    x"7",
        x"5",    x"3",    x"2",    x"0",    x"1",    x"3",    x"4",    x"6",
        x"8",    x"A",    x"C",    x"D",    x"E",    x"C",    x"A",    x"9",
        x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",    x"5",
        x"7",    x"8",    x"A",    x"C",    x"E",    x"E",    x"C",    x"A",
        x"8",    x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",
        x"5",    x"7",    x"9",    x"A",    x"C",    x"E",    x"D",    x"C",
        x"A",    x"8",    x"6",    x"5",    x"6",    x"8",    x"C",    x"C",
        x"8",    x"4",    x"0",    x"4",    x"9",    x"D",    x"B",    x"7",
        x"2",    x"1",    x"6",    x"A",    x"E",    x"A",    x"6",    x"1",
        x"2",    x"7",    x"B",    x"D",    x"9",    x"5",    x"0",    x"3",
        x"8",    x"C",    x"C",    x"8",    x"3",    x"0",    x"5",    x"9",
        x"D",    x"B",    x"7",    x"2",    x"1",    x"6",    x"A",    x"E",
        x"A",    x"6",    x"1",    x"2",    x"7",    x"B",    x"D",    x"9",
        x"4",    x"0",    x"4",    x"8",    x"D",    x"C",    x"8",    x"3",
        x"0",    x"5",    x"9",    x"E",    x"B",    x"6",    x"0",    x"5",
        x"B",    x"C",    x"6",    x"0",    x"5",    x"B",    x"C",    x"6",
        x"0",    x"5",    x"B",    x"C",    x"6",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"F",
        x"F",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",
        x"A",    x"4",    x"1",    x"7",    x"D",    x"A",    x"4",    x"1",
        x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",    x"A",
        x"4",    x"2",    x"C",    x"8",    x"0",    x"9",    x"B",    x"2",
        x"6",    x"E",    x"5",    x"3",    x"C",    x"8",    x"0",    x"9",
        x"B",    x"2",    x"6",    x"F",    x"6",    x"3",    x"C",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"2",    x"B",    x"9",    x"0",    x"8",    x"C",    x"3",
        x"5",    x"E",    x"6",    x"2",    x"B",    x"9",    x"0",    x"8",
        x"C",    x"3",    x"5",    x"E",    x"6",    x"2",    x"B",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"9",    x"0",    x"C",    x"5",    x"6",    x"B",    x"0",
        x"C",    x"5",    x"6",    x"B",    x"1",    x"D",    x"4",    x"7",
        x"A",    x"1",    x"D",    x"4",    x"7",    x"A",    x"2",    x"E",
        x"3",    x"8",    x"9",    x"2",    x"E",    x"3",    x"8",    x"9",
        x"3",    x"E",    x"2",    x"9",    x"8",    x"3",    x"E",    x"2",
        x"9",    x"8",    x"4",    x"D",    x"1",    x"A",    x"7",    x"4",
        x"D",    x"1",    x"A",    x"7",    x"4",    x"C",    x"0",    x"B",
        x"6",    x"1",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"4",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"5",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"4",    x"6",    x"8",    x"9",
        x"B",    x"D",    x"E",    x"D",    x"B",    x"9",    x"7",    x"6",
        x"4",    x"2",    x"0",    x"1",    x"2",    x"4",    x"6",    x"8",
        x"A",    x"B",    x"D",    x"E",    x"C",    x"B",    x"9",    x"7",
        x"5",    x"3",    x"2",    x"0",    x"1",    x"3",    x"4",    x"6",
        x"8",    x"A",    x"C",    x"D",    x"E",    x"C",    x"A",    x"9",
        x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",    x"5",
        x"7",    x"8",    x"A",    x"C",    x"E",    x"E",    x"C",    x"A",
        x"8",    x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",
        x"5",    x"7",    x"9",    x"A",    x"C",    x"E",    x"D",    x"C",
        x"A",    x"8",    x"6",    x"5",    x"6",    x"8",    x"C",    x"C",
        x"8",    x"4",    x"0",    x"4",    x"9",    x"D",    x"B",    x"7",
        x"2",    x"1",    x"6",    x"A",    x"E",    x"A",    x"6",    x"1",
        x"2",    x"7",    x"B",    x"D",    x"9",    x"5",    x"0",    x"3",
        x"8",    x"C",    x"C",    x"8",    x"3",    x"0",    x"5",    x"9",
        x"D",    x"B",    x"7",    x"2",    x"1",    x"6",    x"A",    x"E",
        x"A",    x"6",    x"1",    x"2",    x"7",    x"B",    x"D",    x"9",
        x"4",    x"0",    x"4",    x"8",    x"D",    x"C",    x"8",    x"3",
        x"0",    x"5",    x"9",    x"E",    x"B",    x"6",    x"0",    x"5",
        x"B",    x"C",    x"6",    x"0",    x"5",    x"B",    x"C",    x"6",
        x"0",    x"5",    x"B",    x"C",    x"6",    x"0",    x"1",    x"2",
        x"2",    x"1",    x"0",    x"1",    x"2",    x"2",    x"1",    x"0",
        x"1",    x"2",    x"2",    x"1",    x"0",    x"1",    x"5",    x"C",
        x"C",    x"3",    x"1",    x"2",    x"2",    x"1",    x"0",    x"1",
        x"2",    x"2",    x"1",    x"0",    x"1",    x"2",    x"2",    x"1",
        x"0",    x"1",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",
        x"A",    x"4",    x"1",    x"7",    x"D",    x"A",    x"4",    x"1",
        x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",    x"A",
        x"4",    x"2",    x"C",    x"8",    x"0",    x"9",    x"B",    x"2",
        x"6",    x"E",    x"5",    x"3",    x"C",    x"8",    x"0",    x"9",
        x"B",    x"2",    x"6",    x"F",    x"6",    x"3",    x"C",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"2",    x"B",    x"9",    x"0",    x"8",    x"C",    x"3",
        x"5",    x"E",    x"6",    x"2",    x"B",    x"9",    x"0",    x"8",
        x"C",    x"3",    x"5",    x"E",    x"6",    x"2",    x"B",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"9",    x"0",    x"C",    x"5",    x"6",    x"B",    x"0",
        x"C",    x"5",    x"6",    x"B",    x"1",    x"D",    x"4",    x"7",
        x"A",    x"1",    x"D",    x"4",    x"7",    x"A",    x"2",    x"E",
        x"3",    x"8",    x"9",    x"2",    x"E",    x"3",    x"8",    x"9",
        x"3",    x"E",    x"2",    x"9",    x"8",    x"3",    x"E",    x"2",
        x"9",    x"8",    x"4",    x"D",    x"1",    x"A",    x"7",    x"4",
        x"D",    x"1",    x"A",    x"7",    x"4",    x"C",    x"0",    x"B",
        x"6",    x"1",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"6",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"4",    x"6",    x"8",    x"9",
        x"B",    x"D",    x"E",    x"D",    x"B",    x"9",    x"7",    x"6",
        x"4",    x"2",    x"0",    x"1",    x"2",    x"4",    x"6",    x"8",
        x"A",    x"B",    x"D",    x"E",    x"C",    x"B",    x"9",    x"7",
        x"5",    x"3",    x"2",    x"0",    x"1",    x"3",    x"4",    x"6",
        x"8",    x"A",    x"C",    x"D",    x"E",    x"C",    x"A",    x"9",
        x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",    x"5",
        x"7",    x"8",    x"A",    x"C",    x"E",    x"E",    x"C",    x"A",
        x"8",    x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",
        x"5",    x"7",    x"9",    x"A",    x"C",    x"E",    x"D",    x"C",
        x"A",    x"8",    x"6",    x"5",    x"6",    x"8",    x"C",    x"C",
        x"8",    x"4",    x"0",    x"4",    x"9",    x"D",    x"B",    x"7",
        x"2",    x"1",    x"6",    x"A",    x"E",    x"A",    x"6",    x"1",
        x"2",    x"7",    x"B",    x"D",    x"9",    x"5",    x"0",    x"3",
        x"8",    x"C",    x"C",    x"8",    x"3",    x"0",    x"5",    x"9",
        x"D",    x"B",    x"7",    x"2",    x"1",    x"6",    x"A",    x"E",
        x"A",    x"6",    x"1",    x"2",    x"7",    x"B",    x"D",    x"9",
        x"4",    x"0",    x"4",    x"8",    x"D",    x"C",    x"8",    x"3",
        x"0",    x"5",    x"9",    x"E",    x"B",    x"6",    x"0",    x"5",
        x"B",    x"C",    x"6",    x"0",    x"5",    x"B",    x"C",    x"6",
        x"0",    x"5",    x"B",    x"C",    x"6",    x"0",    x"6",    x"C",
        x"B",    x"5",    x"0",    x"6",    x"C",    x"B",    x"5",    x"0",
        x"6",    x"C",    x"B",    x"5",    x"0",    x"6",    x"C",    x"B",
        x"5",    x"0",    x"6",    x"C",    x"B",    x"5",    x"0",    x"6",
        x"C",    x"B",    x"5",    x"0",    x"6",    x"C",    x"B",    x"5",
        x"1",    x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",
        x"A",    x"4",    x"1",    x"7",    x"D",    x"A",    x"4",    x"1",
        x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",    x"A",
        x"4",    x"2",    x"C",    x"8",    x"0",    x"9",    x"B",    x"2",
        x"6",    x"E",    x"5",    x"3",    x"C",    x"8",    x"0",    x"9",
        x"B",    x"2",    x"6",    x"F",    x"6",    x"3",    x"C",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"2",    x"B",    x"9",    x"0",    x"8",    x"C",    x"3",
        x"5",    x"E",    x"6",    x"2",    x"B",    x"9",    x"0",    x"8",
        x"C",    x"3",    x"5",    x"E",    x"6",    x"2",    x"B",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"9",    x"0",    x"C",    x"5",    x"6",    x"B",    x"0",
        x"C",    x"5",    x"6",    x"B",    x"1",    x"D",    x"4",    x"7",
        x"A",    x"1",    x"D",    x"4",    x"7",    x"A",    x"2",    x"E",
        x"3",    x"8",    x"9",    x"2",    x"E",    x"3",    x"8",    x"9",
        x"3",    x"E",    x"2",    x"9",    x"8",    x"3",    x"E",    x"2",
        x"9",    x"8",    x"4",    x"D",    x"1",    x"A",    x"7",    x"4",
        x"D",    x"1",    x"A",    x"7",    x"4",    x"C",    x"0",    x"B",
        x"6",    x"1",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"1",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"4",    x"6",    x"8",    x"9",
        x"B",    x"D",    x"E",    x"D",    x"B",    x"9",    x"7",    x"6",
        x"4",    x"2",    x"0",    x"1",    x"2",    x"4",    x"6",    x"8",
        x"A",    x"B",    x"D",    x"E",    x"C",    x"B",    x"9",    x"7",
        x"5",    x"3",    x"2",    x"0",    x"1",    x"3",    x"4",    x"6",
        x"8",    x"A",    x"C",    x"D",    x"E",    x"C",    x"A",    x"9",
        x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",    x"5",
        x"7",    x"8",    x"A",    x"C",    x"E",    x"E",    x"C",    x"A",
        x"8",    x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",
        x"5",    x"7",    x"9",    x"A",    x"C",    x"E",    x"D",    x"C",
        x"A",    x"8",    x"6",    x"5",    x"6",    x"8",    x"C",    x"C",
        x"8",    x"4",    x"0",    x"4",    x"9",    x"D",    x"B",    x"7",
        x"2",    x"1",    x"6",    x"A",    x"E",    x"A",    x"6",    x"1",
        x"2",    x"7",    x"B",    x"D",    x"9",    x"5",    x"0",    x"3",
        x"8",    x"C",    x"C",    x"8",    x"3",    x"0",    x"5",    x"9",
        x"D",    x"B",    x"7",    x"2",    x"1",    x"6",    x"A",    x"E",
        x"A",    x"6",    x"1",    x"2",    x"7",    x"B",    x"D",    x"9",
        x"4",    x"0",    x"4",    x"8",    x"D",    x"C",    x"8",    x"3",
        x"0",    x"5",    x"9",    x"E",    x"B",    x"6",    x"0",    x"5",
        x"B",    x"C",    x"6",    x"0",    x"5",    x"B",    x"C",    x"6",
        x"0",    x"5",    x"B",    x"C",    x"6",    x"0",    x"6",    x"C",
        x"B",    x"5",    x"0",    x"6",    x"C",    x"B",    x"5",    x"0",
        x"6",    x"C",    x"B",    x"5",    x"0",    x"6",    x"C",    x"B",
        x"5",    x"0",    x"6",    x"C",    x"B",    x"5",    x"0",    x"6",
        x"C",    x"B",    x"5",    x"0",    x"6",    x"C",    x"B",    x"5",
        x"1",    x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",
        x"A",    x"4",    x"1",    x"7",    x"D",    x"A",    x"4",    x"1",
        x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",    x"A",
        x"4",    x"2",    x"C",    x"8",    x"0",    x"9",    x"B",    x"2",
        x"6",    x"E",    x"5",    x"3",    x"C",    x"8",    x"0",    x"9",
        x"B",    x"2",    x"6",    x"F",    x"6",    x"3",    x"C",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"2",    x"B",    x"9",    x"0",    x"8",    x"C",    x"3",
        x"5",    x"E",    x"6",    x"2",    x"B",    x"9",    x"0",    x"8",
        x"C",    x"3",    x"5",    x"E",    x"6",    x"2",    x"B",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"9",    x"0",    x"C",    x"5",    x"6",    x"B",    x"0",
        x"C",    x"5",    x"6",    x"B",    x"1",    x"D",    x"4",    x"7",
        x"A",    x"1",    x"D",    x"4",    x"7",    x"A",    x"2",    x"E",
        x"3",    x"8",    x"9",    x"2",    x"E",    x"3",    x"8",    x"9",
        x"3",    x"E",    x"2",    x"9",    x"8",    x"3",    x"E",    x"2",
        x"9",    x"8",    x"4",    x"D",    x"1",    x"A",    x"7",    x"4",
        x"D",    x"1",    x"A",    x"7",    x"4",    x"C",    x"0",    x"B",
        x"6",    x"1",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"1",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"4",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"4",    x"6",    x"8",    x"9",
        x"B",    x"D",    x"E",    x"D",    x"B",    x"9",    x"7",    x"6",
        x"4",    x"2",    x"0",    x"1",    x"2",    x"4",    x"6",    x"8",
        x"A",    x"B",    x"D",    x"E",    x"C",    x"B",    x"9",    x"7",
        x"5",    x"3",    x"2",    x"0",    x"1",    x"3",    x"4",    x"6",
        x"8",    x"A",    x"C",    x"D",    x"E",    x"C",    x"A",    x"9",
        x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",    x"5",
        x"7",    x"8",    x"A",    x"C",    x"E",    x"E",    x"C",    x"A",
        x"8",    x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",
        x"5",    x"7",    x"9",    x"A",    x"C",    x"E",    x"D",    x"C",
        x"A",    x"8",    x"6",    x"5",    x"6",    x"8",    x"C",    x"C",
        x"8",    x"4",    x"0",    x"4",    x"9",    x"D",    x"B",    x"7",
        x"2",    x"1",    x"6",    x"A",    x"E",    x"A",    x"6",    x"1",
        x"2",    x"7",    x"B",    x"D",    x"9",    x"5",    x"0",    x"3",
        x"8",    x"C",    x"C",    x"8",    x"3",    x"0",    x"5",    x"9",
        x"D",    x"B",    x"7",    x"2",    x"1",    x"6",    x"A",    x"E",
        x"A",    x"6",    x"1",    x"2",    x"7",    x"B",    x"D",    x"9",
        x"4",    x"0",    x"4",    x"8",    x"D",    x"C",    x"8",    x"3",
        x"0",    x"5",    x"9",    x"E",    x"B",    x"6",    x"0",    x"5",
        x"B",    x"C",    x"6",    x"0",    x"5",    x"B",    x"C",    x"6",
        x"0",    x"5",    x"B",    x"C",    x"6",    x"0",    x"6",    x"C",
        x"B",    x"5",    x"0",    x"6",    x"C",    x"B",    x"5",    x"0",
        x"6",    x"C",    x"B",    x"5",    x"0",    x"6",    x"C",    x"B",
        x"5",    x"0",    x"6",    x"C",    x"B",    x"5",    x"0",    x"6",
        x"C",    x"B",    x"5",    x"0",    x"6",    x"C",    x"B",    x"5",
        x"1",    x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",
        x"A",    x"4",    x"1",    x"7",    x"D",    x"A",    x"4",    x"1",
        x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",    x"A",
        x"4",    x"2",    x"C",    x"8",    x"0",    x"9",    x"B",    x"2",
        x"6",    x"E",    x"5",    x"3",    x"C",    x"8",    x"0",    x"9",
        x"B",    x"2",    x"6",    x"F",    x"6",    x"3",    x"C",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"2",    x"B",    x"9",    x"0",    x"8",    x"C",    x"3",
        x"5",    x"E",    x"6",    x"2",    x"B",    x"9",    x"0",    x"8",
        x"C",    x"3",    x"5",    x"E",    x"6",    x"2",    x"B",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"9",    x"0",    x"C",    x"5",    x"6",    x"B",    x"0",
        x"C",    x"5",    x"6",    x"B",    x"1",    x"D",    x"4",    x"7",
        x"A",    x"1",    x"D",    x"4",    x"7",    x"A",    x"2",    x"E",
        x"3",    x"8",    x"9",    x"2",    x"E",    x"3",    x"8",    x"9",
        x"3",    x"E",    x"2",    x"9",    x"8",    x"3",    x"E",    x"2",
        x"9",    x"8",    x"4",    x"D",    x"1",    x"A",    x"7",    x"4",
        x"D",    x"1",    x"A",    x"7",    x"4",    x"C",    x"0",    x"B",
        x"6",    x"1",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"6",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"4",    x"6",    x"8",    x"9",
        x"B",    x"D",    x"E",    x"D",    x"B",    x"9",    x"7",    x"6",
        x"4",    x"2",    x"0",    x"1",    x"2",    x"4",    x"6",    x"8",
        x"A",    x"B",    x"D",    x"E",    x"C",    x"B",    x"9",    x"7",
        x"5",    x"3",    x"2",    x"0",    x"1",    x"3",    x"4",    x"6",
        x"8",    x"A",    x"C",    x"D",    x"E",    x"C",    x"A",    x"9",
        x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",    x"5",
        x"7",    x"8",    x"A",    x"C",    x"E",    x"E",    x"C",    x"A",
        x"8",    x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",
        x"5",    x"7",    x"9",    x"A",    x"C",    x"E",    x"D",    x"C",
        x"A",    x"8",    x"6",    x"5",    x"6",    x"8",    x"C",    x"C",
        x"8",    x"4",    x"0",    x"4",    x"9",    x"D",    x"B",    x"7",
        x"2",    x"1",    x"6",    x"A",    x"E",    x"A",    x"6",    x"1",
        x"2",    x"7",    x"B",    x"D",    x"9",    x"5",    x"0",    x"3",
        x"8",    x"C",    x"C",    x"8",    x"3",    x"0",    x"5",    x"9",
        x"D",    x"B",    x"7",    x"2",    x"1",    x"6",    x"A",    x"E",
        x"A",    x"6",    x"1",    x"2",    x"7",    x"B",    x"D",    x"9",
        x"4",    x"0",    x"4",    x"8",    x"D",    x"C",    x"8",    x"3",
        x"0",    x"5",    x"9",    x"E",    x"B",    x"6",    x"0",    x"5",
        x"B",    x"C",    x"6",    x"0",    x"5",    x"B",    x"C",    x"6",
        x"0",    x"5",    x"B",    x"C",    x"6",    x"0",    x"6",    x"C",
        x"B",    x"5",    x"0",    x"6",    x"C",    x"B",    x"5",    x"0",
        x"6",    x"C",    x"B",    x"5",    x"0",    x"6",    x"C",    x"B",
        x"5",    x"0",    x"6",    x"C",    x"B",    x"5",    x"0",    x"6",
        x"C",    x"B",    x"5",    x"0",    x"6",    x"C",    x"B",    x"5",
        x"1",    x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",
        x"A",    x"4",    x"1",    x"7",    x"D",    x"A",    x"4",    x"1",
        x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",    x"A",
        x"4",    x"2",    x"C",    x"8",    x"0",    x"9",    x"B",    x"2",
        x"6",    x"E",    x"5",    x"3",    x"C",    x"8",    x"0",    x"9",
        x"B",    x"2",    x"6",    x"F",    x"6",    x"3",    x"C",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"2",    x"B",    x"9",    x"0",    x"8",    x"C",    x"3",
        x"5",    x"E",    x"6",    x"2",    x"B",    x"9",    x"0",    x"8",
        x"C",    x"3",    x"5",    x"E",    x"6",    x"2",    x"B",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"9",    x"0",    x"C",    x"5",    x"6",    x"B",    x"0",
        x"C",    x"5",    x"6",    x"B",    x"1",    x"D",    x"4",    x"7",
        x"A",    x"1",    x"D",    x"4",    x"7",    x"A",    x"2",    x"E",
        x"3",    x"8",    x"9",    x"2",    x"E",    x"3",    x"8",    x"9",
        x"3",    x"E",    x"2",    x"9",    x"8",    x"3",    x"E",    x"2",
        x"9",    x"8",    x"4",    x"D",    x"1",    x"A",    x"7",    x"4",
        x"D",    x"1",    x"A",    x"7",    x"4",    x"C",    x"0",    x"B",
        x"6",    x"1",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"6",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"4",    x"6",    x"8",    x"9",
        x"B",    x"D",    x"E",    x"D",    x"B",    x"9",    x"7",    x"6",
        x"4",    x"2",    x"0",    x"1",    x"2",    x"4",    x"6",    x"8",
        x"A",    x"B",    x"D",    x"E",    x"C",    x"B",    x"9",    x"7",
        x"5",    x"3",    x"2",    x"0",    x"1",    x"3",    x"4",    x"6",
        x"8",    x"A",    x"C",    x"D",    x"E",    x"C",    x"A",    x"9",
        x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",    x"5",
        x"7",    x"8",    x"A",    x"C",    x"E",    x"E",    x"C",    x"A",
        x"8",    x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",
        x"5",    x"7",    x"9",    x"A",    x"C",    x"E",    x"D",    x"C",
        x"A",    x"8",    x"6",    x"5",    x"6",    x"8",    x"C",    x"C",
        x"8",    x"4",    x"0",    x"4",    x"9",    x"D",    x"B",    x"7",
        x"2",    x"1",    x"6",    x"A",    x"E",    x"A",    x"6",    x"1",
        x"2",    x"7",    x"B",    x"D",    x"9",    x"5",    x"0",    x"3",
        x"8",    x"C",    x"C",    x"8",    x"3",    x"0",    x"5",    x"9",
        x"D",    x"B",    x"7",    x"2",    x"1",    x"6",    x"A",    x"E",
        x"A",    x"6",    x"1",    x"2",    x"7",    x"B",    x"D",    x"9",
        x"4",    x"0",    x"4",    x"8",    x"D",    x"C",    x"8",    x"3",
        x"0",    x"5",    x"9",    x"E",    x"B",    x"6",    x"0",    x"5",
        x"B",    x"C",    x"6",    x"0",    x"5",    x"B",    x"C",    x"6",
        x"0",    x"5",    x"B",    x"C",    x"6",    x"0",    x"6",    x"C",
        x"B",    x"5",    x"0",    x"6",    x"C",    x"B",    x"5",    x"0",
        x"6",    x"C",    x"B",    x"5",    x"0",    x"6",    x"C",    x"B",
        x"5",    x"0",    x"6",    x"C",    x"B",    x"5",    x"0",    x"6",
        x"C",    x"B",    x"5",    x"0",    x"6",    x"C",    x"B",    x"5",
        x"1",    x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",
        x"A",    x"4",    x"1",    x"7",    x"D",    x"A",    x"4",    x"1",
        x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",    x"A",
        x"4",    x"2",    x"C",    x"8",    x"0",    x"9",    x"B",    x"2",
        x"6",    x"E",    x"5",    x"3",    x"C",    x"8",    x"0",    x"9",
        x"B",    x"2",    x"6",    x"F",    x"6",    x"3",    x"C",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"2",    x"B",    x"9",    x"0",    x"8",    x"C",    x"3",
        x"5",    x"E",    x"6",    x"2",    x"B",    x"9",    x"0",    x"8",
        x"C",    x"3",    x"5",    x"E",    x"6",    x"2",    x"B",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"9",    x"0",    x"C",    x"5",    x"6",    x"B",    x"0",
        x"C",    x"5",    x"6",    x"B",    x"1",    x"D",    x"4",    x"7",
        x"A",    x"1",    x"D",    x"4",    x"7",    x"A",    x"2",    x"E",
        x"3",    x"8",    x"9",    x"2",    x"E",    x"3",    x"8",    x"9",
        x"3",    x"E",    x"2",    x"9",    x"8",    x"3",    x"E",    x"2",
        x"9",    x"8",    x"4",    x"D",    x"1",    x"A",    x"7",    x"4",
        x"D",    x"1",    x"A",    x"7",    x"4",    x"C",    x"0",    x"B",
        x"6",    x"1",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"3",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"4",    x"6",    x"8",    x"9",
        x"B",    x"D",    x"E",    x"D",    x"B",    x"9",    x"7",    x"6",
        x"4",    x"2",    x"0",    x"1",    x"2",    x"4",    x"6",    x"8",
        x"A",    x"B",    x"D",    x"E",    x"C",    x"B",    x"9",    x"7",
        x"5",    x"3",    x"2",    x"0",    x"1",    x"3",    x"4",    x"6",
        x"8",    x"A",    x"C",    x"D",    x"E",    x"C",    x"A",    x"9",
        x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",    x"5",
        x"7",    x"8",    x"A",    x"C",    x"E",    x"E",    x"C",    x"A",
        x"8",    x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",
        x"5",    x"7",    x"9",    x"A",    x"C",    x"E",    x"D",    x"C",
        x"A",    x"8",    x"6",    x"5",    x"6",    x"8",    x"C",    x"C",
        x"8",    x"4",    x"0",    x"4",    x"9",    x"D",    x"B",    x"7",
        x"2",    x"1",    x"6",    x"A",    x"E",    x"A",    x"6",    x"1",
        x"2",    x"7",    x"B",    x"D",    x"9",    x"5",    x"0",    x"3",
        x"8",    x"C",    x"C",    x"8",    x"3",    x"0",    x"5",    x"9",
        x"D",    x"B",    x"7",    x"2",    x"1",    x"6",    x"A",    x"E",
        x"A",    x"6",    x"1",    x"2",    x"7",    x"B",    x"D",    x"9",
        x"4",    x"0",    x"4",    x"8",    x"D",    x"C",    x"8",    x"3",
        x"0",    x"5",    x"9",    x"E",    x"B",    x"6",    x"0",    x"5",
        x"B",    x"C",    x"6",    x"0",    x"5",    x"B",    x"C",    x"6",
        x"0",    x"5",    x"B",    x"C",    x"6",    x"0",    x"6",    x"C",
        x"B",    x"5",    x"0",    x"6",    x"C",    x"B",    x"5",    x"0",
        x"6",    x"C",    x"B",    x"5",    x"0",    x"6",    x"C",    x"B",
        x"5",    x"0",    x"6",    x"C",    x"B",    x"5",    x"0",    x"6",
        x"C",    x"B",    x"5",    x"0",    x"6",    x"C",    x"B",    x"5",
        x"1",    x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",
        x"A",    x"4",    x"1",    x"7",    x"D",    x"A",    x"4",    x"1",
        x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",    x"A",
        x"4",    x"2",    x"C",    x"8",    x"0",    x"9",    x"B",    x"2",
        x"6",    x"E",    x"5",    x"3",    x"C",    x"8",    x"0",    x"9",
        x"B",    x"2",    x"6",    x"F",    x"6",    x"3",    x"C",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"2",    x"B",    x"9",    x"0",    x"8",    x"C",    x"3",
        x"5",    x"E",    x"6",    x"2",    x"B",    x"9",    x"0",    x"8",
        x"C",    x"3",    x"5",    x"E",    x"6",    x"2",    x"B",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"9",    x"0",    x"C",    x"5",    x"6",    x"B",    x"0",
        x"C",    x"5",    x"6",    x"B",    x"1",    x"D",    x"4",    x"7",
        x"A",    x"1",    x"D",    x"4",    x"7",    x"A",    x"2",    x"E",
        x"3",    x"8",    x"9",    x"2",    x"E",    x"3",    x"8",    x"9",
        x"3",    x"E",    x"2",    x"9",    x"8",    x"3",    x"E",    x"2",
        x"9",    x"8",    x"4",    x"D",    x"1",    x"A",    x"7",    x"4",
        x"D",    x"1",    x"A",    x"7",    x"4",    x"C",    x"0",    x"B",
        x"6",    x"1",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"3",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"5",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"4",    x"6",    x"8",    x"9",
        x"B",    x"D",    x"E",    x"D",    x"B",    x"9",    x"7",    x"6",
        x"4",    x"2",    x"0",    x"1",    x"2",    x"4",    x"6",    x"8",
        x"A",    x"B",    x"D",    x"E",    x"C",    x"B",    x"9",    x"7",
        x"5",    x"3",    x"2",    x"0",    x"1",    x"3",    x"4",    x"6",
        x"8",    x"A",    x"C",    x"D",    x"E",    x"C",    x"A",    x"9",
        x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",    x"5",
        x"7",    x"8",    x"A",    x"C",    x"E",    x"E",    x"C",    x"A",
        x"8",    x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",
        x"5",    x"7",    x"9",    x"A",    x"C",    x"E",    x"D",    x"C",
        x"A",    x"8",    x"6",    x"5",    x"6",    x"8",    x"C",    x"C",
        x"8",    x"4",    x"0",    x"4",    x"9",    x"D",    x"B",    x"7",
        x"2",    x"1",    x"6",    x"A",    x"E",    x"A",    x"6",    x"1",
        x"2",    x"7",    x"B",    x"D",    x"9",    x"5",    x"0",    x"3",
        x"8",    x"C",    x"C",    x"8",    x"3",    x"0",    x"5",    x"9",
        x"D",    x"B",    x"7",    x"2",    x"1",    x"6",    x"A",    x"E",
        x"A",    x"6",    x"1",    x"2",    x"7",    x"B",    x"D",    x"9",
        x"4",    x"0",    x"4",    x"8",    x"D",    x"C",    x"8",    x"3",
        x"0",    x"5",    x"9",    x"E",    x"B",    x"6",    x"0",    x"5",
        x"B",    x"C",    x"6",    x"0",    x"5",    x"B",    x"C",    x"6",
        x"0",    x"5",    x"B",    x"C",    x"6",    x"0",    x"6",    x"C",
        x"B",    x"5",    x"0",    x"6",    x"C",    x"B",    x"5",    x"0",
        x"6",    x"C",    x"B",    x"5",    x"0",    x"6",    x"C",    x"B",
        x"5",    x"0",    x"6",    x"C",    x"B",    x"5",    x"0",    x"6",
        x"C",    x"B",    x"5",    x"0",    x"6",    x"C",    x"B",    x"5",
        x"1",    x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",
        x"A",    x"4",    x"1",    x"7",    x"D",    x"A",    x"4",    x"1",
        x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",    x"A",
        x"4",    x"2",    x"C",    x"8",    x"0",    x"9",    x"B",    x"2",
        x"6",    x"E",    x"5",    x"3",    x"C",    x"8",    x"0",    x"9",
        x"B",    x"2",    x"6",    x"F",    x"6",    x"3",    x"C",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"2",    x"B",    x"9",    x"0",    x"8",    x"C",    x"3",
        x"5",    x"E",    x"6",    x"2",    x"B",    x"9",    x"0",    x"8",
        x"C",    x"3",    x"5",    x"E",    x"6",    x"2",    x"B",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"9",    x"0",    x"C",    x"5",    x"6",    x"B",    x"0",
        x"C",    x"5",    x"6",    x"B",    x"1",    x"D",    x"4",    x"7",
        x"A",    x"1",    x"D",    x"4",    x"7",    x"A",    x"2",    x"E",
        x"3",    x"8",    x"9",    x"2",    x"E",    x"3",    x"8",    x"9",
        x"3",    x"E",    x"2",    x"9",    x"8",    x"3",    x"E",    x"2",
        x"9",    x"8",    x"4",    x"D",    x"1",    x"A",    x"7",    x"4",
        x"D",    x"1",    x"A",    x"7",    x"4",    x"C",    x"0",    x"B",
        x"6",    x"1",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"5",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"4",    x"6",    x"8",    x"9",
        x"B",    x"D",    x"E",    x"D",    x"B",    x"9",    x"7",    x"6",
        x"4",    x"2",    x"0",    x"1",    x"2",    x"4",    x"6",    x"8",
        x"A",    x"B",    x"D",    x"E",    x"C",    x"B",    x"9",    x"7",
        x"5",    x"3",    x"2",    x"0",    x"1",    x"3",    x"4",    x"6",
        x"8",    x"A",    x"C",    x"D",    x"E",    x"C",    x"A",    x"9",
        x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",    x"5",
        x"7",    x"8",    x"A",    x"C",    x"E",    x"E",    x"C",    x"A",
        x"8",    x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",
        x"5",    x"7",    x"9",    x"A",    x"C",    x"E",    x"D",    x"C",
        x"A",    x"8",    x"6",    x"5",    x"6",    x"8",    x"C",    x"C",
        x"8",    x"4",    x"0",    x"4",    x"9",    x"D",    x"B",    x"7",
        x"2",    x"1",    x"6",    x"A",    x"E",    x"A",    x"6",    x"1",
        x"2",    x"7",    x"B",    x"D",    x"9",    x"5",    x"0",    x"3",
        x"8",    x"C",    x"C",    x"8",    x"3",    x"0",    x"5",    x"9",
        x"D",    x"B",    x"7",    x"2",    x"1",    x"6",    x"A",    x"E",
        x"A",    x"6",    x"1",    x"2",    x"7",    x"B",    x"D",    x"9",
        x"4",    x"0",    x"4",    x"8",    x"D",    x"C",    x"8",    x"3",
        x"0",    x"5",    x"9",    x"E",    x"B",    x"6",    x"0",    x"5",
        x"B",    x"C",    x"6",    x"0",    x"5",    x"B",    x"C",    x"6",
        x"0",    x"5",    x"B",    x"C",    x"6",    x"0",    x"6",    x"C",
        x"B",    x"5",    x"0",    x"6",    x"C",    x"B",    x"5",    x"0",
        x"6",    x"C",    x"B",    x"5",    x"0",    x"6",    x"C",    x"B",
        x"5",    x"0",    x"6",    x"C",    x"B",    x"5",    x"0",    x"6",
        x"C",    x"B",    x"5",    x"0",    x"6",    x"C",    x"B",    x"5",
        x"1",    x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",
        x"A",    x"4",    x"1",    x"7",    x"D",    x"A",    x"4",    x"1",
        x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",    x"A",
        x"4",    x"2",    x"C",    x"8",    x"0",    x"9",    x"B",    x"2",
        x"6",    x"E",    x"5",    x"3",    x"C",    x"8",    x"0",    x"9",
        x"B",    x"2",    x"6",    x"F",    x"6",    x"3",    x"C",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"2",    x"B",    x"9",    x"0",    x"8",    x"C",    x"3",
        x"5",    x"E",    x"6",    x"2",    x"B",    x"9",    x"0",    x"8",
        x"C",    x"3",    x"5",    x"E",    x"6",    x"2",    x"B",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"9",    x"0",    x"C",    x"5",    x"6",    x"B",    x"0",
        x"C",    x"5",    x"6",    x"B",    x"1",    x"D",    x"4",    x"7",
        x"A",    x"1",    x"D",    x"4",    x"7",    x"A",    x"2",    x"E",
        x"3",    x"8",    x"9",    x"2",    x"E",    x"3",    x"8",    x"9",
        x"3",    x"E",    x"2",    x"9",    x"8",    x"3",    x"E",    x"2",
        x"9",    x"8",    x"4",    x"D",    x"1",    x"A",    x"7",    x"4",
        x"D",    x"1",    x"A",    x"7",    x"4",    x"C",    x"0",    x"B",
        x"6",    x"1",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"1",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"4",    x"6",    x"8",    x"9",
        x"B",    x"D",    x"E",    x"D",    x"B",    x"9",    x"7",    x"6",
        x"4",    x"2",    x"0",    x"1",    x"2",    x"4",    x"6",    x"8",
        x"A",    x"B",    x"D",    x"E",    x"C",    x"B",    x"9",    x"7",
        x"5",    x"3",    x"2",    x"0",    x"1",    x"3",    x"4",    x"6",
        x"8",    x"A",    x"C",    x"D",    x"E",    x"C",    x"A",    x"9",
        x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",    x"5",
        x"7",    x"8",    x"A",    x"C",    x"E",    x"E",    x"C",    x"A",
        x"8",    x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",
        x"5",    x"7",    x"9",    x"A",    x"C",    x"E",    x"D",    x"C",
        x"A",    x"8",    x"6",    x"5",    x"6",    x"8",    x"C",    x"C",
        x"8",    x"4",    x"0",    x"4",    x"9",    x"D",    x"B",    x"7",
        x"2",    x"1",    x"6",    x"A",    x"E",    x"A",    x"6",    x"1",
        x"2",    x"7",    x"B",    x"D",    x"9",    x"5",    x"0",    x"3",
        x"8",    x"C",    x"C",    x"8",    x"3",    x"0",    x"5",    x"9",
        x"D",    x"B",    x"7",    x"2",    x"1",    x"6",    x"A",    x"E",
        x"A",    x"6",    x"1",    x"2",    x"7",    x"B",    x"D",    x"9",
        x"4",    x"0",    x"4",    x"8",    x"D",    x"C",    x"8",    x"3",
        x"0",    x"5",    x"9",    x"E",    x"B",    x"6",    x"0",    x"5",
        x"B",    x"C",    x"6",    x"0",    x"5",    x"B",    x"C",    x"6",
        x"0",    x"5",    x"B",    x"C",    x"6",    x"0",    x"6",    x"C",
        x"B",    x"5",    x"0",    x"6",    x"C",    x"B",    x"5",    x"0",
        x"6",    x"C",    x"B",    x"5",    x"0",    x"6",    x"C",    x"B",
        x"5",    x"0",    x"6",    x"C",    x"B",    x"5",    x"0",    x"6",
        x"C",    x"B",    x"5",    x"0",    x"6",    x"C",    x"B",    x"5",
        x"1",    x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",
        x"A",    x"4",    x"1",    x"7",    x"D",    x"A",    x"4",    x"1",
        x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",    x"A",
        x"4",    x"2",    x"C",    x"8",    x"0",    x"9",    x"B",    x"2",
        x"6",    x"E",    x"5",    x"3",    x"C",    x"8",    x"0",    x"9",
        x"B",    x"2",    x"6",    x"F",    x"6",    x"3",    x"C",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"2",    x"B",    x"9",    x"0",    x"8",    x"C",    x"3",
        x"5",    x"E",    x"6",    x"2",    x"B",    x"9",    x"0",    x"8",
        x"C",    x"3",    x"5",    x"E",    x"6",    x"2",    x"B",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"9",    x"0",    x"C",    x"5",    x"6",    x"B",    x"0",
        x"C",    x"5",    x"6",    x"B",    x"1",    x"D",    x"4",    x"7",
        x"A",    x"1",    x"D",    x"4",    x"7",    x"A",    x"2",    x"E",
        x"3",    x"8",    x"9",    x"2",    x"E",    x"3",    x"8",    x"9",
        x"3",    x"E",    x"2",    x"9",    x"8",    x"3",    x"E",    x"2",
        x"9",    x"8",    x"4",    x"D",    x"1",    x"A",    x"7",    x"4",
        x"D",    x"1",    x"A",    x"7",    x"4",    x"C",    x"0",    x"B",
        x"6",    x"1",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"1",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"5",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"4",    x"6",    x"8",    x"9",
        x"B",    x"D",    x"E",    x"D",    x"B",    x"9",    x"7",    x"6",
        x"4",    x"2",    x"0",    x"1",    x"2",    x"4",    x"6",    x"8",
        x"A",    x"B",    x"D",    x"E",    x"C",    x"B",    x"9",    x"7",
        x"5",    x"3",    x"2",    x"0",    x"1",    x"3",    x"4",    x"6",
        x"8",    x"A",    x"C",    x"D",    x"E",    x"C",    x"A",    x"9",
        x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",    x"5",
        x"7",    x"8",    x"A",    x"C",    x"E",    x"E",    x"C",    x"A",
        x"8",    x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",
        x"5",    x"7",    x"9",    x"A",    x"C",    x"E",    x"D",    x"C",
        x"A",    x"8",    x"6",    x"5",    x"6",    x"8",    x"C",    x"C",
        x"8",    x"4",    x"0",    x"4",    x"9",    x"D",    x"B",    x"7",
        x"2",    x"1",    x"6",    x"A",    x"E",    x"A",    x"6",    x"1",
        x"2",    x"7",    x"B",    x"D",    x"9",    x"5",    x"0",    x"3",
        x"8",    x"C",    x"C",    x"8",    x"3",    x"0",    x"5",    x"9",
        x"D",    x"B",    x"7",    x"2",    x"1",    x"6",    x"A",    x"E",
        x"A",    x"6",    x"1",    x"2",    x"7",    x"B",    x"D",    x"9",
        x"4",    x"0",    x"4",    x"8",    x"D",    x"C",    x"8",    x"3",
        x"0",    x"5",    x"9",    x"E",    x"B",    x"6",    x"0",    x"5",
        x"B",    x"C",    x"6",    x"0",    x"5",    x"B",    x"C",    x"6",
        x"0",    x"5",    x"B",    x"C",    x"6",    x"0",    x"6",    x"C",
        x"B",    x"5",    x"0",    x"6",    x"C",    x"B",    x"5",    x"0",
        x"6",    x"C",    x"B",    x"5",    x"0",    x"6",    x"C",    x"B",
        x"5",    x"0",    x"6",    x"C",    x"B",    x"5",    x"0",    x"6",
        x"C",    x"B",    x"5",    x"0",    x"6",    x"C",    x"B",    x"5",
        x"1",    x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",
        x"A",    x"4",    x"1",    x"7",    x"D",    x"A",    x"4",    x"1",
        x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",    x"A",
        x"4",    x"2",    x"C",    x"8",    x"0",    x"9",    x"B",    x"2",
        x"6",    x"E",    x"5",    x"3",    x"C",    x"8",    x"0",    x"9",
        x"B",    x"2",    x"6",    x"F",    x"6",    x"3",    x"C",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"2",    x"B",    x"9",    x"0",    x"8",    x"C",    x"3",
        x"5",    x"E",    x"6",    x"2",    x"B",    x"9",    x"0",    x"8",
        x"C",    x"3",    x"5",    x"E",    x"6",    x"2",    x"B",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"9",    x"0",    x"C",    x"5",    x"6",    x"B",    x"0",
        x"C",    x"5",    x"6",    x"B",    x"1",    x"D",    x"4",    x"7",
        x"A",    x"1",    x"D",    x"4",    x"7",    x"A",    x"2",    x"E",
        x"3",    x"8",    x"9",    x"2",    x"E",    x"3",    x"8",    x"9",
        x"3",    x"E",    x"2",    x"9",    x"8",    x"3",    x"E",    x"2",
        x"9",    x"8",    x"4",    x"D",    x"1",    x"A",    x"7",    x"4",
        x"D",    x"1",    x"A",    x"7",    x"4",    x"C",    x"0",    x"B",
        x"6",    x"1",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"5",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"4",    x"6",    x"8",    x"9",
        x"B",    x"D",    x"E",    x"D",    x"B",    x"9",    x"7",    x"6",
        x"4",    x"2",    x"0",    x"1",    x"2",    x"4",    x"6",    x"8",
        x"A",    x"B",    x"D",    x"E",    x"C",    x"B",    x"9",    x"7",
        x"5",    x"3",    x"2",    x"0",    x"1",    x"3",    x"4",    x"6",
        x"8",    x"A",    x"C",    x"D",    x"E",    x"C",    x"A",    x"9",
        x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",    x"5",
        x"7",    x"8",    x"A",    x"C",    x"E",    x"E",    x"C",    x"A",
        x"8",    x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",
        x"5",    x"7",    x"9",    x"A",    x"C",    x"E",    x"D",    x"C",
        x"A",    x"8",    x"6",    x"5",    x"6",    x"8",    x"C",    x"C",
        x"8",    x"4",    x"0",    x"4",    x"9",    x"D",    x"B",    x"7",
        x"2",    x"1",    x"6",    x"A",    x"E",    x"A",    x"6",    x"1",
        x"2",    x"7",    x"B",    x"D",    x"9",    x"5",    x"0",    x"3",
        x"8",    x"C",    x"C",    x"8",    x"3",    x"0",    x"5",    x"9",
        x"D",    x"B",    x"7",    x"2",    x"1",    x"6",    x"A",    x"E",
        x"A",    x"6",    x"1",    x"2",    x"7",    x"B",    x"D",    x"9",
        x"4",    x"0",    x"4",    x"8",    x"D",    x"C",    x"8",    x"3",
        x"0",    x"5",    x"9",    x"E",    x"B",    x"6",    x"0",    x"5",
        x"B",    x"C",    x"6",    x"0",    x"5",    x"B",    x"C",    x"6",
        x"0",    x"5",    x"B",    x"C",    x"6",    x"0",    x"6",    x"C",
        x"B",    x"5",    x"0",    x"6",    x"C",    x"B",    x"5",    x"0",
        x"6",    x"C",    x"B",    x"5",    x"0",    x"6",    x"C",    x"B",
        x"5",    x"0",    x"6",    x"C",    x"B",    x"5",    x"0",    x"6",
        x"C",    x"B",    x"5",    x"0",    x"6",    x"C",    x"B",    x"5",
        x"1",    x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",
        x"A",    x"4",    x"1",    x"7",    x"D",    x"A",    x"4",    x"1",
        x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",    x"A",
        x"4",    x"2",    x"C",    x"8",    x"0",    x"9",    x"B",    x"2",
        x"6",    x"E",    x"5",    x"3",    x"C",    x"8",    x"0",    x"9",
        x"B",    x"2",    x"6",    x"F",    x"6",    x"3",    x"C",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"2",    x"B",    x"9",    x"0",    x"8",    x"C",    x"3",
        x"5",    x"E",    x"6",    x"2",    x"B",    x"9",    x"0",    x"8",
        x"C",    x"3",    x"5",    x"E",    x"6",    x"2",    x"B",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"9",    x"0",    x"C",    x"5",    x"6",    x"B",    x"0",
        x"C",    x"5",    x"6",    x"B",    x"1",    x"D",    x"4",    x"7",
        x"A",    x"1",    x"D",    x"4",    x"7",    x"A",    x"2",    x"E",
        x"3",    x"8",    x"9",    x"2",    x"E",    x"3",    x"8",    x"9",
        x"3",    x"E",    x"2",    x"9",    x"8",    x"3",    x"E",    x"2",
        x"9",    x"8",    x"4",    x"D",    x"1",    x"A",    x"7",    x"4",
        x"D",    x"1",    x"A",    x"7",    x"4",    x"C",    x"0",    x"B",
        x"6",    x"1",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"1",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"4",    x"6",    x"8",    x"9",
        x"B",    x"D",    x"E",    x"D",    x"B",    x"9",    x"7",    x"6",
        x"4",    x"2",    x"0",    x"1",    x"2",    x"4",    x"6",    x"8",
        x"A",    x"B",    x"D",    x"E",    x"C",    x"B",    x"9",    x"7",
        x"5",    x"3",    x"2",    x"0",    x"1",    x"3",    x"4",    x"6",
        x"8",    x"A",    x"C",    x"D",    x"E",    x"C",    x"A",    x"9",
        x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",    x"5",
        x"7",    x"8",    x"A",    x"C",    x"E",    x"E",    x"C",    x"A",
        x"8",    x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",
        x"5",    x"7",    x"9",    x"A",    x"C",    x"E",    x"D",    x"C",
        x"A",    x"8",    x"6",    x"5",    x"6",    x"8",    x"C",    x"C",
        x"8",    x"4",    x"0",    x"4",    x"9",    x"D",    x"B",    x"7",
        x"2",    x"1",    x"6",    x"A",    x"E",    x"A",    x"6",    x"1",
        x"2",    x"7",    x"B",    x"D",    x"9",    x"5",    x"0",    x"3",
        x"8",    x"C",    x"C",    x"8",    x"3",    x"0",    x"5",    x"9",
        x"D",    x"B",    x"7",    x"2",    x"1",    x"6",    x"A",    x"E",
        x"A",    x"6",    x"1",    x"2",    x"7",    x"B",    x"D",    x"9",
        x"4",    x"0",    x"4",    x"8",    x"D",    x"C",    x"8",    x"3",
        x"0",    x"5",    x"9",    x"E",    x"B",    x"6",    x"0",    x"5",
        x"B",    x"C",    x"6",    x"0",    x"5",    x"B",    x"C",    x"6",
        x"0",    x"5",    x"B",    x"C",    x"6",    x"0",    x"6",    x"C",
        x"B",    x"5",    x"0",    x"6",    x"C",    x"B",    x"5",    x"0",
        x"6",    x"C",    x"B",    x"5",    x"0",    x"6",    x"C",    x"B",
        x"5",    x"0",    x"6",    x"C",    x"B",    x"5",    x"0",    x"6",
        x"C",    x"B",    x"5",    x"0",    x"6",    x"C",    x"B",    x"5",
        x"1",    x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",
        x"A",    x"4",    x"1",    x"7",    x"D",    x"A",    x"4",    x"1",
        x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",    x"A",
        x"4",    x"2",    x"C",    x"8",    x"0",    x"9",    x"B",    x"2",
        x"6",    x"E",    x"5",    x"3",    x"C",    x"8",    x"0",    x"9",
        x"B",    x"2",    x"6",    x"F",    x"6",    x"3",    x"C",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"2",    x"B",    x"9",    x"0",    x"8",    x"C",    x"3",
        x"5",    x"E",    x"6",    x"2",    x"B",    x"9",    x"0",    x"8",
        x"C",    x"3",    x"5",    x"E",    x"6",    x"2",    x"B",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"9",    x"0",    x"C",    x"5",    x"6",    x"B",    x"0",
        x"C",    x"5",    x"6",    x"B",    x"1",    x"D",    x"4",    x"7",
        x"A",    x"1",    x"D",    x"4",    x"7",    x"A",    x"2",    x"E",
        x"3",    x"8",    x"9",    x"2",    x"E",    x"3",    x"8",    x"9",
        x"3",    x"E",    x"2",    x"9",    x"8",    x"3",    x"E",    x"2",
        x"9",    x"8",    x"4",    x"D",    x"1",    x"A",    x"7",    x"4",
        x"D",    x"1",    x"A",    x"7",    x"4",    x"C",    x"0",    x"B",
        x"6",    x"1",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"1",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"5",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"4",    x"6",    x"8",    x"9",
        x"B",    x"D",    x"E",    x"D",    x"B",    x"9",    x"7",    x"6",
        x"4",    x"2",    x"0",    x"1",    x"2",    x"4",    x"6",    x"8",
        x"A",    x"B",    x"D",    x"E",    x"C",    x"B",    x"9",    x"7",
        x"5",    x"3",    x"2",    x"0",    x"1",    x"3",    x"4",    x"6",
        x"8",    x"A",    x"C",    x"D",    x"E",    x"C",    x"A",    x"9",
        x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",    x"5",
        x"7",    x"8",    x"A",    x"C",    x"E",    x"E",    x"C",    x"A",
        x"8",    x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",
        x"5",    x"7",    x"9",    x"A",    x"C",    x"E",    x"D",    x"C",
        x"A",    x"8",    x"6",    x"5",    x"6",    x"8",    x"C",    x"C",
        x"8",    x"4",    x"0",    x"4",    x"9",    x"D",    x"B",    x"7",
        x"2",    x"1",    x"6",    x"A",    x"E",    x"A",    x"6",    x"1",
        x"2",    x"7",    x"B",    x"D",    x"9",    x"5",    x"0",    x"3",
        x"8",    x"C",    x"C",    x"8",    x"3",    x"0",    x"5",    x"9",
        x"D",    x"B",    x"7",    x"2",    x"1",    x"6",    x"A",    x"E",
        x"A",    x"6",    x"1",    x"2",    x"7",    x"B",    x"D",    x"9",
        x"4",    x"0",    x"4",    x"8",    x"D",    x"C",    x"8",    x"3",
        x"0",    x"5",    x"9",    x"E",    x"B",    x"6",    x"0",    x"5",
        x"B",    x"C",    x"6",    x"0",    x"5",    x"B",    x"C",    x"6",
        x"0",    x"5",    x"B",    x"C",    x"6",    x"0",    x"6",    x"C",
        x"B",    x"5",    x"0",    x"6",    x"C",    x"B",    x"5",    x"0",
        x"6",    x"C",    x"B",    x"5",    x"0",    x"6",    x"C",    x"B",
        x"5",    x"0",    x"6",    x"C",    x"B",    x"5",    x"0",    x"6",
        x"C",    x"B",    x"5",    x"0",    x"6",    x"C",    x"B",    x"5",
        x"1",    x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",
        x"A",    x"4",    x"1",    x"7",    x"D",    x"A",    x"4",    x"1",
        x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",    x"A",
        x"4",    x"2",    x"C",    x"8",    x"0",    x"9",    x"B",    x"2",
        x"6",    x"E",    x"5",    x"3",    x"C",    x"8",    x"0",    x"9",
        x"B",    x"2",    x"6",    x"F",    x"6",    x"3",    x"C",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"2",    x"B",    x"9",    x"0",    x"8",    x"C",    x"3",
        x"5",    x"E",    x"6",    x"2",    x"B",    x"9",    x"0",    x"8",
        x"C",    x"3",    x"5",    x"E",    x"6",    x"2",    x"B",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"9",    x"0",    x"C",    x"5",    x"6",    x"B",    x"0",
        x"C",    x"5",    x"6",    x"B",    x"1",    x"D",    x"4",    x"7",
        x"A",    x"1",    x"D",    x"4",    x"7",    x"A",    x"2",    x"E",
        x"3",    x"8",    x"9",    x"2",    x"E",    x"3",    x"8",    x"9",
        x"3",    x"E",    x"2",    x"9",    x"8",    x"3",    x"E",    x"2",
        x"9",    x"8",    x"4",    x"D",    x"1",    x"A",    x"7",    x"4",
        x"D",    x"1",    x"A",    x"7",    x"4",    x"C",    x"0",    x"B",
        x"6",    x"1",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"5",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"4",    x"6",    x"8",    x"9",
        x"B",    x"D",    x"E",    x"D",    x"B",    x"9",    x"7",    x"6",
        x"4",    x"2",    x"0",    x"1",    x"2",    x"4",    x"6",    x"8",
        x"A",    x"B",    x"D",    x"E",    x"C",    x"B",    x"9",    x"7",
        x"5",    x"3",    x"2",    x"0",    x"1",    x"3",    x"4",    x"6",
        x"8",    x"A",    x"C",    x"D",    x"E",    x"C",    x"A",    x"9",
        x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",    x"5",
        x"7",    x"8",    x"A",    x"C",    x"E",    x"E",    x"C",    x"A",
        x"8",    x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",
        x"5",    x"7",    x"9",    x"A",    x"C",    x"E",    x"D",    x"C",
        x"A",    x"8",    x"6",    x"5",    x"6",    x"8",    x"C",    x"C",
        x"8",    x"4",    x"0",    x"4",    x"9",    x"D",    x"B",    x"7",
        x"2",    x"1",    x"6",    x"A",    x"E",    x"A",    x"6",    x"1",
        x"2",    x"7",    x"B",    x"D",    x"9",    x"5",    x"0",    x"3",
        x"8",    x"C",    x"C",    x"8",    x"3",    x"0",    x"5",    x"9",
        x"D",    x"B",    x"7",    x"2",    x"1",    x"6",    x"A",    x"E",
        x"A",    x"6",    x"1",    x"2",    x"7",    x"B",    x"D",    x"9",
        x"4",    x"0",    x"4",    x"8",    x"D",    x"C",    x"8",    x"3",
        x"0",    x"5",    x"9",    x"E",    x"B",    x"6",    x"0",    x"5",
        x"B",    x"C",    x"6",    x"0",    x"5",    x"B",    x"C",    x"6",
        x"0",    x"5",    x"B",    x"C",    x"6",    x"0",    x"6",    x"C",
        x"B",    x"5",    x"0",    x"6",    x"C",    x"B",    x"5",    x"0",
        x"6",    x"C",    x"B",    x"5",    x"0",    x"6",    x"C",    x"B",
        x"5",    x"0",    x"6",    x"C",    x"B",    x"5",    x"0",    x"6",
        x"C",    x"B",    x"5",    x"0",    x"6",    x"C",    x"B",    x"5",
        x"1",    x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",
        x"A",    x"4",    x"1",    x"7",    x"D",    x"A",    x"4",    x"1",
        x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",    x"A",
        x"4",    x"2",    x"C",    x"8",    x"0",    x"9",    x"B",    x"2",
        x"6",    x"E",    x"5",    x"3",    x"C",    x"8",    x"0",    x"9",
        x"B",    x"2",    x"6",    x"F",    x"6",    x"3",    x"C",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"2",    x"B",    x"9",    x"0",    x"8",    x"C",    x"3",
        x"5",    x"E",    x"6",    x"2",    x"B",    x"9",    x"0",    x"8",
        x"C",    x"3",    x"5",    x"E",    x"6",    x"2",    x"B",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"9",    x"0",    x"C",    x"5",    x"6",    x"B",    x"0",
        x"C",    x"5",    x"6",    x"B",    x"1",    x"D",    x"4",    x"7",
        x"A",    x"1",    x"D",    x"4",    x"7",    x"A",    x"2",    x"E",
        x"3",    x"8",    x"9",    x"2",    x"E",    x"3",    x"8",    x"9",
        x"3",    x"E",    x"2",    x"9",    x"8",    x"3",    x"E",    x"2",
        x"9",    x"8",    x"4",    x"D",    x"1",    x"A",    x"7",    x"4",
        x"D",    x"1",    x"A",    x"7",    x"4",    x"C",    x"0",    x"B",
        x"6",    x"1",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"1",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"4",    x"6",    x"8",    x"9",
        x"B",    x"D",    x"E",    x"D",    x"B",    x"9",    x"7",    x"6",
        x"4",    x"2",    x"0",    x"1",    x"2",    x"4",    x"6",    x"8",
        x"A",    x"B",    x"D",    x"E",    x"C",    x"B",    x"9",    x"7",
        x"5",    x"3",    x"2",    x"0",    x"1",    x"3",    x"4",    x"6",
        x"8",    x"A",    x"C",    x"D",    x"E",    x"C",    x"A",    x"9",
        x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",    x"5",
        x"7",    x"8",    x"A",    x"C",    x"E",    x"E",    x"C",    x"A",
        x"8",    x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",
        x"5",    x"7",    x"9",    x"A",    x"C",    x"E",    x"D",    x"C",
        x"A",    x"8",    x"6",    x"5",    x"6",    x"8",    x"C",    x"C",
        x"8",    x"4",    x"0",    x"4",    x"9",    x"D",    x"B",    x"7",
        x"2",    x"1",    x"6",    x"A",    x"E",    x"A",    x"6",    x"1",
        x"2",    x"7",    x"B",    x"D",    x"9",    x"5",    x"0",    x"3",
        x"8",    x"C",    x"C",    x"8",    x"3",    x"0",    x"5",    x"9",
        x"D",    x"B",    x"7",    x"2",    x"1",    x"6",    x"A",    x"E",
        x"A",    x"6",    x"1",    x"2",    x"7",    x"B",    x"D",    x"9",
        x"4",    x"0",    x"4",    x"8",    x"D",    x"C",    x"8",    x"3",
        x"0",    x"5",    x"9",    x"E",    x"B",    x"6",    x"0",    x"5",
        x"B",    x"C",    x"6",    x"0",    x"5",    x"B",    x"C",    x"6",
        x"0",    x"5",    x"B",    x"C",    x"6",    x"0",    x"6",    x"C",
        x"B",    x"5",    x"0",    x"6",    x"C",    x"B",    x"5",    x"0",
        x"6",    x"C",    x"B",    x"5",    x"0",    x"6",    x"C",    x"B",
        x"5",    x"0",    x"6",    x"C",    x"B",    x"5",    x"0",    x"6",
        x"C",    x"B",    x"5",    x"0",    x"6",    x"C",    x"B",    x"5",
        x"1",    x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",
        x"A",    x"4",    x"1",    x"7",    x"D",    x"A",    x"4",    x"1",
        x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",    x"A",
        x"4",    x"2",    x"C",    x"8",    x"0",    x"9",    x"B",    x"2",
        x"6",    x"E",    x"5",    x"3",    x"C",    x"8",    x"0",    x"9",
        x"B",    x"2",    x"6",    x"F",    x"6",    x"3",    x"C",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"2",    x"B",    x"9",    x"0",    x"8",    x"C",    x"3",
        x"5",    x"E",    x"6",    x"2",    x"B",    x"9",    x"0",    x"8",
        x"C",    x"3",    x"5",    x"E",    x"6",    x"2",    x"B",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"9",    x"0",    x"C",    x"5",    x"6",    x"B",    x"0",
        x"C",    x"5",    x"6",    x"B",    x"1",    x"D",    x"4",    x"7",
        x"A",    x"1",    x"D",    x"4",    x"7",    x"A",    x"2",    x"E",
        x"3",    x"8",    x"9",    x"2",    x"E",    x"3",    x"8",    x"9",
        x"3",    x"E",    x"2",    x"9",    x"8",    x"3",    x"E",    x"2",
        x"9",    x"8",    x"4",    x"D",    x"1",    x"A",    x"7",    x"4",
        x"D",    x"1",    x"A",    x"7",    x"4",    x"C",    x"0",    x"B",
        x"6",    x"1",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"1",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"5",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"4",    x"6",    x"8",    x"9",
        x"B",    x"D",    x"E",    x"D",    x"B",    x"9",    x"7",    x"6",
        x"4",    x"2",    x"0",    x"1",    x"2",    x"4",    x"6",    x"8",
        x"A",    x"B",    x"D",    x"E",    x"C",    x"B",    x"9",    x"7",
        x"5",    x"3",    x"2",    x"0",    x"1",    x"3",    x"4",    x"6",
        x"8",    x"A",    x"C",    x"D",    x"E",    x"C",    x"A",    x"9",
        x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",    x"5",
        x"7",    x"8",    x"A",    x"C",    x"E",    x"E",    x"C",    x"A",
        x"8",    x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",
        x"5",    x"7",    x"9",    x"A",    x"C",    x"E",    x"D",    x"C",
        x"A",    x"8",    x"6",    x"5",    x"6",    x"8",    x"C",    x"C",
        x"8",    x"4",    x"0",    x"4",    x"9",    x"D",    x"B",    x"7",
        x"2",    x"1",    x"6",    x"A",    x"E",    x"A",    x"6",    x"1",
        x"2",    x"7",    x"B",    x"D",    x"9",    x"5",    x"0",    x"3",
        x"8",    x"C",    x"C",    x"8",    x"3",    x"0",    x"5",    x"9",
        x"D",    x"B",    x"7",    x"2",    x"1",    x"6",    x"A",    x"E",
        x"A",    x"6",    x"1",    x"2",    x"7",    x"B",    x"D",    x"9",
        x"4",    x"0",    x"4",    x"8",    x"D",    x"C",    x"8",    x"3",
        x"0",    x"5",    x"9",    x"E",    x"B",    x"6",    x"0",    x"5",
        x"B",    x"C",    x"6",    x"0",    x"5",    x"B",    x"C",    x"6",
        x"0",    x"5",    x"B",    x"C",    x"6",    x"0",    x"6",    x"C",
        x"B",    x"5",    x"0",    x"6",    x"C",    x"B",    x"5",    x"0",
        x"6",    x"C",    x"B",    x"5",    x"0",    x"6",    x"C",    x"B",
        x"5",    x"0",    x"6",    x"C",    x"B",    x"5",    x"0",    x"6",
        x"C",    x"B",    x"5",    x"0",    x"6",    x"C",    x"B",    x"5",
        x"1",    x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",
        x"A",    x"4",    x"1",    x"7",    x"D",    x"A",    x"4",    x"1",
        x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",    x"A",
        x"4",    x"2",    x"C",    x"8",    x"0",    x"9",    x"B",    x"2",
        x"6",    x"E",    x"5",    x"3",    x"C",    x"8",    x"0",    x"9",
        x"B",    x"2",    x"6",    x"F",    x"6",    x"3",    x"C",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"2",    x"B",    x"9",    x"0",    x"8",    x"C",    x"3",
        x"5",    x"E",    x"6",    x"2",    x"B",    x"9",    x"0",    x"8",
        x"C",    x"3",    x"5",    x"E",    x"6",    x"2",    x"B",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"9",    x"0",    x"C",    x"5",    x"6",    x"B",    x"0",
        x"C",    x"5",    x"6",    x"B",    x"1",    x"D",    x"4",    x"7",
        x"A",    x"1",    x"D",    x"4",    x"7",    x"A",    x"2",    x"E",
        x"3",    x"8",    x"9",    x"2",    x"E",    x"3",    x"8",    x"9",
        x"3",    x"E",    x"2",    x"9",    x"8",    x"3",    x"E",    x"2",
        x"9",    x"8",    x"4",    x"D",    x"1",    x"A",    x"7",    x"4",
        x"D",    x"1",    x"A",    x"7",    x"4",    x"C",    x"0",    x"B",
        x"6",    x"1",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"5",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"4",    x"6",    x"8",    x"9",
        x"B",    x"D",    x"E",    x"D",    x"B",    x"9",    x"7",    x"6",
        x"4",    x"2",    x"0",    x"1",    x"2",    x"4",    x"6",    x"8",
        x"A",    x"B",    x"D",    x"E",    x"C",    x"B",    x"9",    x"7",
        x"5",    x"3",    x"2",    x"0",    x"1",    x"3",    x"4",    x"6",
        x"8",    x"A",    x"C",    x"D",    x"E",    x"C",    x"A",    x"9",
        x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",    x"5",
        x"7",    x"8",    x"A",    x"C",    x"E",    x"E",    x"C",    x"A",
        x"8",    x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",
        x"5",    x"7",    x"9",    x"A",    x"C",    x"E",    x"D",    x"C",
        x"A",    x"8",    x"6",    x"5",    x"6",    x"8",    x"C",    x"C",
        x"8",    x"4",    x"0",    x"4",    x"9",    x"D",    x"B",    x"7",
        x"2",    x"1",    x"6",    x"A",    x"E",    x"A",    x"6",    x"1",
        x"2",    x"7",    x"B",    x"D",    x"9",    x"5",    x"0",    x"3",
        x"8",    x"C",    x"C",    x"8",    x"3",    x"0",    x"5",    x"9",
        x"D",    x"B",    x"7",    x"2",    x"1",    x"6",    x"A",    x"E",
        x"A",    x"6",    x"1",    x"2",    x"7",    x"B",    x"D",    x"9",
        x"4",    x"0",    x"4",    x"8",    x"D",    x"C",    x"8",    x"3",
        x"0",    x"5",    x"9",    x"E",    x"B",    x"6",    x"0",    x"5",
        x"B",    x"C",    x"6",    x"0",    x"5",    x"B",    x"C",    x"6",
        x"0",    x"5",    x"B",    x"C",    x"6",    x"0",    x"6",    x"C",
        x"B",    x"5",    x"0",    x"6",    x"C",    x"B",    x"5",    x"0",
        x"6",    x"C",    x"B",    x"5",    x"0",    x"6",    x"C",    x"B",
        x"5",    x"0",    x"6",    x"C",    x"B",    x"5",    x"0",    x"6",
        x"C",    x"B",    x"5",    x"0",    x"6",    x"C",    x"B",    x"5",
        x"1",    x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",
        x"A",    x"4",    x"1",    x"7",    x"D",    x"A",    x"4",    x"1",
        x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",    x"A",
        x"4",    x"2",    x"C",    x"8",    x"0",    x"9",    x"B",    x"2",
        x"6",    x"E",    x"5",    x"3",    x"C",    x"8",    x"0",    x"9",
        x"B",    x"2",    x"6",    x"F",    x"6",    x"3",    x"C",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"2",    x"B",    x"9",    x"0",    x"8",    x"C",    x"3",
        x"5",    x"E",    x"6",    x"2",    x"B",    x"9",    x"0",    x"8",
        x"C",    x"3",    x"5",    x"E",    x"6",    x"2",    x"B",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"9",    x"0",    x"C",    x"5",    x"6",    x"B",    x"0",
        x"C",    x"5",    x"6",    x"B",    x"1",    x"D",    x"4",    x"7",
        x"A",    x"1",    x"D",    x"4",    x"7",    x"A",    x"2",    x"E",
        x"3",    x"8",    x"9",    x"2",    x"E",    x"3",    x"8",    x"9",
        x"3",    x"E",    x"2",    x"9",    x"8",    x"3",    x"E",    x"2",
        x"9",    x"8",    x"4",    x"D",    x"1",    x"A",    x"7",    x"4",
        x"D",    x"1",    x"A",    x"7",    x"4",    x"C",    x"0",    x"B",
        x"6",    x"1",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"2",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"4",    x"6",    x"8",    x"9",
        x"B",    x"D",    x"E",    x"D",    x"B",    x"9",    x"7",    x"6",
        x"4",    x"2",    x"0",    x"1",    x"2",    x"4",    x"6",    x"8",
        x"A",    x"B",    x"D",    x"E",    x"C",    x"B",    x"9",    x"7",
        x"5",    x"3",    x"2",    x"0",    x"1",    x"3",    x"4",    x"6",
        x"8",    x"A",    x"C",    x"D",    x"E",    x"C",    x"A",    x"9",
        x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",    x"5",
        x"7",    x"8",    x"A",    x"C",    x"E",    x"E",    x"C",    x"A",
        x"8",    x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",
        x"5",    x"7",    x"9",    x"A",    x"C",    x"E",    x"D",    x"C",
        x"A",    x"8",    x"6",    x"5",    x"6",    x"8",    x"C",    x"C",
        x"8",    x"4",    x"0",    x"4",    x"9",    x"D",    x"B",    x"7",
        x"2",    x"1",    x"6",    x"A",    x"E",    x"A",    x"6",    x"1",
        x"2",    x"7",    x"B",    x"D",    x"9",    x"5",    x"0",    x"3",
        x"8",    x"C",    x"C",    x"8",    x"3",    x"0",    x"5",    x"9",
        x"D",    x"B",    x"7",    x"2",    x"1",    x"6",    x"A",    x"E",
        x"A",    x"6",    x"1",    x"2",    x"7",    x"B",    x"D",    x"9",
        x"4",    x"0",    x"4",    x"8",    x"D",    x"C",    x"8",    x"3",
        x"0",    x"5",    x"9",    x"E",    x"B",    x"6",    x"0",    x"5",
        x"B",    x"C",    x"6",    x"0",    x"5",    x"B",    x"C",    x"6",
        x"0",    x"5",    x"B",    x"C",    x"6",    x"0",    x"6",    x"C",
        x"B",    x"5",    x"0",    x"6",    x"C",    x"B",    x"5",    x"0",
        x"6",    x"C",    x"B",    x"5",    x"0",    x"6",    x"C",    x"B",
        x"5",    x"0",    x"6",    x"C",    x"B",    x"5",    x"0",    x"6",
        x"C",    x"B",    x"5",    x"0",    x"6",    x"C",    x"B",    x"5",
        x"1",    x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",
        x"A",    x"4",    x"1",    x"7",    x"D",    x"A",    x"4",    x"1",
        x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",    x"A",
        x"4",    x"2",    x"C",    x"8",    x"0",    x"9",    x"B",    x"2",
        x"6",    x"E",    x"5",    x"3",    x"C",    x"8",    x"0",    x"9",
        x"B",    x"2",    x"6",    x"F",    x"6",    x"3",    x"C",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"2",    x"B",    x"9",    x"0",    x"8",    x"C",    x"3",
        x"5",    x"E",    x"6",    x"2",    x"B",    x"9",    x"0",    x"8",
        x"C",    x"3",    x"5",    x"E",    x"6",    x"2",    x"B",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"9",    x"0",    x"C",    x"5",    x"6",    x"B",    x"0",
        x"C",    x"5",    x"6",    x"B",    x"1",    x"D",    x"4",    x"7",
        x"A",    x"1",    x"D",    x"4",    x"7",    x"A",    x"2",    x"E",
        x"3",    x"8",    x"9",    x"2",    x"E",    x"3",    x"8",    x"9",
        x"3",    x"E",    x"2",    x"9",    x"8",    x"3",    x"E",    x"2",
        x"9",    x"8",    x"4",    x"D",    x"1",    x"A",    x"7",    x"4",
        x"D",    x"1",    x"A",    x"7",    x"4",    x"C",    x"0",    x"B",
        x"6",    x"1",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"5",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"4",    x"6",    x"8",    x"9",
        x"B",    x"D",    x"E",    x"D",    x"B",    x"9",    x"7",    x"6",
        x"4",    x"2",    x"0",    x"1",    x"2",    x"4",    x"6",    x"8",
        x"A",    x"B",    x"D",    x"E",    x"C",    x"B",    x"9",    x"7",
        x"5",    x"3",    x"2",    x"0",    x"1",    x"3",    x"4",    x"6",
        x"8",    x"A",    x"C",    x"D",    x"E",    x"C",    x"A",    x"9",
        x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",    x"5",
        x"7",    x"8",    x"A",    x"C",    x"E",    x"E",    x"C",    x"A",
        x"8",    x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",
        x"5",    x"7",    x"9",    x"A",    x"C",    x"E",    x"D",    x"C",
        x"A",    x"8",    x"6",    x"5",    x"6",    x"8",    x"C",    x"C",
        x"8",    x"4",    x"0",    x"4",    x"9",    x"D",    x"B",    x"7",
        x"2",    x"1",    x"6",    x"A",    x"E",    x"A",    x"6",    x"1",
        x"2",    x"7",    x"B",    x"D",    x"9",    x"5",    x"0",    x"3",
        x"8",    x"C",    x"C",    x"8",    x"3",    x"0",    x"5",    x"9",
        x"D",    x"B",    x"7",    x"2",    x"1",    x"6",    x"A",    x"E",
        x"A",    x"6",    x"1",    x"2",    x"7",    x"B",    x"D",    x"9",
        x"4",    x"0",    x"4",    x"8",    x"D",    x"C",    x"8",    x"3",
        x"0",    x"5",    x"9",    x"E",    x"B",    x"6",    x"0",    x"5",
        x"B",    x"C",    x"6",    x"0",    x"5",    x"B",    x"C",    x"6",
        x"0",    x"5",    x"B",    x"C",    x"6",    x"0",    x"6",    x"C",
        x"B",    x"5",    x"0",    x"6",    x"C",    x"B",    x"5",    x"0",
        x"6",    x"C",    x"B",    x"5",    x"0",    x"6",    x"C",    x"B",
        x"5",    x"0",    x"6",    x"C",    x"B",    x"5",    x"0",    x"6",
        x"C",    x"B",    x"5",    x"0",    x"6",    x"C",    x"B",    x"5",
        x"1",    x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",
        x"A",    x"4",    x"1",    x"7",    x"D",    x"A",    x"4",    x"1",
        x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",    x"A",
        x"4",    x"2",    x"C",    x"8",    x"0",    x"9",    x"B",    x"2",
        x"6",    x"E",    x"5",    x"3",    x"C",    x"8",    x"0",    x"9",
        x"B",    x"2",    x"6",    x"F",    x"6",    x"3",    x"C",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"2",    x"B",    x"9",    x"0",    x"8",    x"C",    x"3",
        x"5",    x"E",    x"6",    x"2",    x"B",    x"9",    x"0",    x"8",
        x"C",    x"3",    x"5",    x"E",    x"6",    x"2",    x"B",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"9",    x"0",    x"C",    x"5",    x"6",    x"B",    x"0",
        x"C",    x"5",    x"6",    x"B",    x"1",    x"D",    x"4",    x"7",
        x"A",    x"1",    x"D",    x"4",    x"7",    x"A",    x"2",    x"E",
        x"3",    x"8",    x"9",    x"2",    x"E",    x"3",    x"8",    x"9",
        x"3",    x"E",    x"2",    x"9",    x"8",    x"3",    x"E",    x"2",
        x"9",    x"8",    x"4",    x"D",    x"1",    x"A",    x"7",    x"4",
        x"D",    x"1",    x"A",    x"7",    x"4",    x"C",    x"0",    x"B",
        x"6",    x"1",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"5",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"4",    x"6",    x"8",    x"9",
        x"B",    x"D",    x"E",    x"D",    x"B",    x"9",    x"7",    x"6",
        x"4",    x"2",    x"0",    x"1",    x"2",    x"4",    x"6",    x"8",
        x"A",    x"B",    x"D",    x"E",    x"C",    x"B",    x"9",    x"7",
        x"5",    x"3",    x"2",    x"0",    x"1",    x"3",    x"4",    x"6",
        x"8",    x"A",    x"C",    x"D",    x"E",    x"C",    x"A",    x"9",
        x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",    x"5",
        x"7",    x"8",    x"A",    x"C",    x"E",    x"E",    x"C",    x"A",
        x"8",    x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",
        x"5",    x"7",    x"9",    x"A",    x"C",    x"E",    x"D",    x"C",
        x"A",    x"8",    x"6",    x"5",    x"6",    x"8",    x"C",    x"C",
        x"8",    x"4",    x"0",    x"4",    x"9",    x"D",    x"B",    x"7",
        x"2",    x"1",    x"6",    x"A",    x"E",    x"A",    x"6",    x"1",
        x"2",    x"7",    x"B",    x"D",    x"9",    x"5",    x"0",    x"3",
        x"8",    x"C",    x"C",    x"8",    x"3",    x"0",    x"5",    x"9",
        x"D",    x"B",    x"7",    x"2",    x"1",    x"6",    x"A",    x"E",
        x"A",    x"6",    x"1",    x"2",    x"7",    x"B",    x"D",    x"9",
        x"4",    x"0",    x"4",    x"8",    x"D",    x"C",    x"8",    x"3",
        x"0",    x"5",    x"9",    x"E",    x"B",    x"6",    x"0",    x"5",
        x"B",    x"C",    x"6",    x"0",    x"5",    x"B",    x"C",    x"6",
        x"0",    x"5",    x"B",    x"C",    x"6",    x"0",    x"6",    x"C",
        x"B",    x"5",    x"0",    x"6",    x"C",    x"B",    x"5",    x"0",
        x"6",    x"C",    x"B",    x"5",    x"0",    x"6",    x"C",    x"B",
        x"5",    x"0",    x"6",    x"C",    x"B",    x"5",    x"0",    x"6",
        x"C",    x"B",    x"5",    x"0",    x"6",    x"C",    x"B",    x"5",
        x"1",    x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",
        x"A",    x"4",    x"1",    x"7",    x"D",    x"A",    x"4",    x"1",
        x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",    x"A",
        x"4",    x"2",    x"C",    x"8",    x"0",    x"9",    x"B",    x"2",
        x"6",    x"E",    x"5",    x"3",    x"C",    x"8",    x"0",    x"9",
        x"B",    x"2",    x"6",    x"F",    x"6",    x"3",    x"C",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"2",    x"B",    x"9",    x"0",    x"8",    x"C",    x"3",
        x"5",    x"E",    x"6",    x"2",    x"B",    x"9",    x"0",    x"8",
        x"C",    x"3",    x"5",    x"E",    x"6",    x"2",    x"B",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"9",    x"0",    x"C",    x"5",    x"6",    x"B",    x"0",
        x"C",    x"5",    x"6",    x"B",    x"1",    x"D",    x"4",    x"7",
        x"A",    x"1",    x"D",    x"4",    x"7",    x"A",    x"2",    x"E",
        x"3",    x"8",    x"9",    x"2",    x"E",    x"3",    x"8",    x"9",
        x"3",    x"E",    x"2",    x"9",    x"8",    x"3",    x"E",    x"2",
        x"9",    x"8",    x"4",    x"D",    x"1",    x"A",    x"7",    x"4",
        x"D",    x"1",    x"A",    x"7",    x"4",    x"C",    x"0",    x"B",
        x"6",    x"1",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"3",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"4",    x"6",    x"8",    x"9",
        x"B",    x"D",    x"E",    x"D",    x"B",    x"9",    x"7",    x"6",
        x"4",    x"2",    x"0",    x"1",    x"2",    x"4",    x"6",    x"8",
        x"A",    x"B",    x"D",    x"E",    x"C",    x"B",    x"9",    x"7",
        x"5",    x"3",    x"2",    x"0",    x"1",    x"3",    x"4",    x"6",
        x"8",    x"A",    x"C",    x"D",    x"E",    x"C",    x"A",    x"9",
        x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",    x"5",
        x"7",    x"8",    x"A",    x"C",    x"E",    x"E",    x"C",    x"A",
        x"8",    x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",
        x"5",    x"7",    x"9",    x"A",    x"C",    x"E",    x"D",    x"C",
        x"A",    x"8",    x"6",    x"5",    x"6",    x"8",    x"C",    x"C",
        x"8",    x"4",    x"0",    x"4",    x"9",    x"D",    x"B",    x"7",
        x"2",    x"1",    x"6",    x"A",    x"E",    x"A",    x"6",    x"1",
        x"2",    x"7",    x"B",    x"D",    x"9",    x"5",    x"0",    x"3",
        x"8",    x"C",    x"C",    x"8",    x"3",    x"0",    x"5",    x"9",
        x"D",    x"B",    x"7",    x"2",    x"1",    x"6",    x"A",    x"E",
        x"A",    x"6",    x"1",    x"2",    x"7",    x"B",    x"D",    x"9",
        x"4",    x"0",    x"4",    x"8",    x"D",    x"C",    x"8",    x"3",
        x"0",    x"5",    x"9",    x"E",    x"B",    x"6",    x"0",    x"5",
        x"B",    x"C",    x"6",    x"0",    x"5",    x"B",    x"C",    x"6",
        x"0",    x"5",    x"B",    x"C",    x"6",    x"0",    x"6",    x"C",
        x"B",    x"5",    x"0",    x"6",    x"C",    x"B",    x"5",    x"0",
        x"6",    x"C",    x"B",    x"5",    x"0",    x"6",    x"C",    x"B",
        x"5",    x"0",    x"6",    x"C",    x"B",    x"5",    x"0",    x"6",
        x"C",    x"B",    x"5",    x"0",    x"6",    x"C",    x"B",    x"5",
        x"1",    x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",
        x"A",    x"4",    x"1",    x"7",    x"D",    x"A",    x"4",    x"1",
        x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",    x"A",
        x"4",    x"2",    x"C",    x"8",    x"0",    x"9",    x"B",    x"2",
        x"6",    x"E",    x"5",    x"3",    x"C",    x"8",    x"0",    x"9",
        x"B",    x"2",    x"6",    x"F",    x"6",    x"3",    x"C",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"2",    x"B",    x"9",    x"0",    x"8",    x"C",    x"3",
        x"5",    x"E",    x"6",    x"2",    x"B",    x"9",    x"0",    x"8",
        x"C",    x"3",    x"5",    x"E",    x"6",    x"2",    x"B",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"9",    x"0",    x"C",    x"5",    x"6",    x"B",    x"0",
        x"C",    x"5",    x"6",    x"B",    x"1",    x"D",    x"4",    x"7",
        x"A",    x"1",    x"D",    x"4",    x"7",    x"A",    x"2",    x"E",
        x"3",    x"8",    x"9",    x"2",    x"E",    x"3",    x"8",    x"9",
        x"3",    x"E",    x"2",    x"9",    x"8",    x"3",    x"E",    x"2",
        x"9",    x"8",    x"4",    x"D",    x"1",    x"A",    x"7",    x"4",
        x"D",    x"1",    x"A",    x"7",    x"4",    x"C",    x"0",    x"B",
        x"6",    x"1",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"3",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"6",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"4",    x"6",    x"8",    x"9",
        x"B",    x"D",    x"E",    x"D",    x"B",    x"9",    x"7",    x"6",
        x"4",    x"2",    x"0",    x"1",    x"2",    x"4",    x"6",    x"8",
        x"A",    x"B",    x"D",    x"E",    x"C",    x"B",    x"9",    x"7",
        x"5",    x"3",    x"2",    x"0",    x"1",    x"3",    x"4",    x"6",
        x"8",    x"A",    x"C",    x"D",    x"E",    x"C",    x"A",    x"9",
        x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",    x"5",
        x"7",    x"8",    x"A",    x"C",    x"E",    x"E",    x"C",    x"A",
        x"8",    x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",
        x"5",    x"7",    x"9",    x"A",    x"C",    x"E",    x"D",    x"C",
        x"A",    x"8",    x"6",    x"5",    x"6",    x"8",    x"C",    x"C",
        x"8",    x"4",    x"0",    x"4",    x"9",    x"D",    x"B",    x"7",
        x"2",    x"1",    x"6",    x"A",    x"E",    x"A",    x"6",    x"1",
        x"2",    x"7",    x"B",    x"D",    x"9",    x"5",    x"0",    x"3",
        x"8",    x"C",    x"C",    x"8",    x"3",    x"0",    x"5",    x"9",
        x"D",    x"B",    x"7",    x"2",    x"1",    x"6",    x"A",    x"E",
        x"A",    x"6",    x"1",    x"2",    x"7",    x"B",    x"D",    x"9",
        x"4",    x"0",    x"4",    x"8",    x"D",    x"C",    x"8",    x"3",
        x"0",    x"5",    x"9",    x"E",    x"B",    x"6",    x"0",    x"5",
        x"B",    x"C",    x"6",    x"0",    x"5",    x"B",    x"C",    x"6",
        x"0",    x"5",    x"B",    x"C",    x"6",    x"0",    x"6",    x"C",
        x"B",    x"5",    x"0",    x"6",    x"C",    x"B",    x"5",    x"0",
        x"6",    x"C",    x"B",    x"5",    x"0",    x"6",    x"C",    x"B",
        x"5",    x"0",    x"6",    x"C",    x"B",    x"5",    x"0",    x"6",
        x"C",    x"B",    x"5",    x"0",    x"6",    x"C",    x"B",    x"5",
        x"1",    x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",
        x"A",    x"4",    x"1",    x"7",    x"D",    x"A",    x"4",    x"1",
        x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",    x"A",
        x"4",    x"2",    x"C",    x"8",    x"0",    x"9",    x"B",    x"2",
        x"6",    x"E",    x"5",    x"3",    x"C",    x"8",    x"0",    x"9",
        x"B",    x"2",    x"6",    x"F",    x"6",    x"3",    x"C",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"2",    x"B",    x"9",    x"0",    x"8",    x"C",    x"3",
        x"5",    x"E",    x"6",    x"2",    x"B",    x"9",    x"0",    x"8",
        x"C",    x"3",    x"5",    x"E",    x"6",    x"2",    x"B",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"9",    x"0",    x"C",    x"5",    x"6",    x"B",    x"0",
        x"C",    x"5",    x"6",    x"B",    x"1",    x"D",    x"4",    x"7",
        x"A",    x"1",    x"D",    x"4",    x"7",    x"A",    x"2",    x"E",
        x"3",    x"8",    x"9",    x"2",    x"E",    x"3",    x"8",    x"9",
        x"3",    x"E",    x"2",    x"9",    x"8",    x"3",    x"E",    x"2",
        x"9",    x"8",    x"4",    x"D",    x"1",    x"A",    x"7",    x"4",
        x"D",    x"1",    x"A",    x"7",    x"4",    x"C",    x"0",    x"B",
        x"6",    x"1",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"6",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"1",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"4",    x"6",    x"8",    x"9",
        x"B",    x"D",    x"E",    x"D",    x"B",    x"9",    x"7",    x"6",
        x"4",    x"2",    x"0",    x"1",    x"2",    x"4",    x"6",    x"8",
        x"A",    x"B",    x"D",    x"E",    x"C",    x"B",    x"9",    x"7",
        x"5",    x"3",    x"2",    x"0",    x"1",    x"3",    x"4",    x"6",
        x"8",    x"A",    x"C",    x"D",    x"E",    x"C",    x"A",    x"9",
        x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",    x"5",
        x"7",    x"8",    x"A",    x"C",    x"E",    x"E",    x"C",    x"A",
        x"8",    x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",
        x"5",    x"7",    x"9",    x"A",    x"C",    x"E",    x"D",    x"C",
        x"A",    x"8",    x"6",    x"5",    x"6",    x"8",    x"C",    x"C",
        x"8",    x"4",    x"0",    x"4",    x"9",    x"D",    x"B",    x"7",
        x"2",    x"1",    x"6",    x"A",    x"E",    x"A",    x"6",    x"1",
        x"2",    x"7",    x"B",    x"D",    x"9",    x"5",    x"0",    x"3",
        x"8",    x"C",    x"C",    x"8",    x"3",    x"0",    x"5",    x"9",
        x"D",    x"B",    x"7",    x"2",    x"1",    x"6",    x"A",    x"E",
        x"A",    x"6",    x"1",    x"2",    x"7",    x"B",    x"D",    x"9",
        x"4",    x"0",    x"4",    x"8",    x"D",    x"C",    x"8",    x"3",
        x"0",    x"5",    x"9",    x"E",    x"B",    x"6",    x"0",    x"5",
        x"B",    x"C",    x"6",    x"0",    x"5",    x"B",    x"C",    x"6",
        x"0",    x"5",    x"B",    x"C",    x"6",    x"0",    x"6",    x"C",
        x"B",    x"5",    x"0",    x"6",    x"C",    x"B",    x"5",    x"0",
        x"6",    x"C",    x"B",    x"5",    x"0",    x"6",    x"C",    x"B",
        x"5",    x"0",    x"6",    x"C",    x"B",    x"5",    x"0",    x"6",
        x"C",    x"B",    x"5",    x"0",    x"6",    x"C",    x"B",    x"5",
        x"1",    x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",
        x"A",    x"4",    x"1",    x"7",    x"D",    x"A",    x"4",    x"1",
        x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",    x"A",
        x"4",    x"2",    x"C",    x"8",    x"0",    x"9",    x"B",    x"2",
        x"6",    x"E",    x"5",    x"3",    x"C",    x"8",    x"0",    x"9",
        x"B",    x"2",    x"6",    x"F",    x"6",    x"3",    x"C",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"2",    x"B",    x"9",    x"0",    x"8",    x"C",    x"3",
        x"5",    x"E",    x"6",    x"2",    x"B",    x"9",    x"0",    x"8",
        x"C",    x"3",    x"5",    x"E",    x"6",    x"2",    x"B",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"9",    x"0",    x"C",    x"5",    x"6",    x"B",    x"0",
        x"C",    x"5",    x"6",    x"B",    x"1",    x"D",    x"4",    x"7",
        x"A",    x"1",    x"D",    x"4",    x"7",    x"A",    x"2",    x"E",
        x"3",    x"8",    x"9",    x"2",    x"E",    x"3",    x"8",    x"9",
        x"3",    x"E",    x"2",    x"9",    x"8",    x"3",    x"E",    x"2",
        x"9",    x"8",    x"4",    x"D",    x"1",    x"A",    x"7",    x"4",
        x"D",    x"1",    x"A",    x"7",    x"4",    x"C",    x"0",    x"B",
        x"6",    x"1",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"1",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"5",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"4",    x"6",    x"8",    x"9",
        x"B",    x"D",    x"E",    x"D",    x"B",    x"9",    x"7",    x"6",
        x"4",    x"2",    x"0",    x"1",    x"2",    x"4",    x"6",    x"8",
        x"A",    x"B",    x"D",    x"E",    x"C",    x"B",    x"9",    x"7",
        x"5",    x"3",    x"2",    x"0",    x"1",    x"3",    x"4",    x"6",
        x"8",    x"A",    x"C",    x"D",    x"E",    x"C",    x"A",    x"9",
        x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",    x"5",
        x"7",    x"8",    x"A",    x"C",    x"E",    x"E",    x"C",    x"A",
        x"8",    x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",
        x"5",    x"7",    x"9",    x"A",    x"C",    x"E",    x"D",    x"C",
        x"A",    x"8",    x"6",    x"5",    x"6",    x"8",    x"C",    x"C",
        x"8",    x"4",    x"0",    x"4",    x"9",    x"D",    x"B",    x"7",
        x"2",    x"1",    x"6",    x"A",    x"E",    x"A",    x"6",    x"1",
        x"2",    x"7",    x"B",    x"D",    x"9",    x"5",    x"0",    x"3",
        x"8",    x"C",    x"C",    x"8",    x"3",    x"0",    x"5",    x"9",
        x"D",    x"B",    x"7",    x"2",    x"1",    x"6",    x"A",    x"E",
        x"A",    x"6",    x"1",    x"2",    x"7",    x"B",    x"D",    x"9",
        x"4",    x"0",    x"4",    x"8",    x"D",    x"C",    x"8",    x"3",
        x"0",    x"5",    x"9",    x"E",    x"B",    x"6",    x"0",    x"5",
        x"B",    x"C",    x"6",    x"0",    x"5",    x"B",    x"C",    x"6",
        x"0",    x"5",    x"B",    x"C",    x"6",    x"0",    x"6",    x"C",
        x"B",    x"5",    x"0",    x"6",    x"C",    x"B",    x"5",    x"0",
        x"6",    x"C",    x"B",    x"5",    x"0",    x"6",    x"C",    x"B",
        x"5",    x"0",    x"6",    x"C",    x"B",    x"5",    x"0",    x"6",
        x"C",    x"B",    x"5",    x"0",    x"6",    x"C",    x"B",    x"5",
        x"1",    x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",
        x"A",    x"4",    x"1",    x"7",    x"D",    x"A",    x"4",    x"1",
        x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",    x"A",
        x"4",    x"2",    x"C",    x"8",    x"0",    x"9",    x"B",    x"2",
        x"6",    x"E",    x"5",    x"3",    x"C",    x"8",    x"0",    x"9",
        x"B",    x"2",    x"6",    x"F",    x"6",    x"3",    x"C",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"2",    x"B",    x"9",    x"0",    x"8",    x"C",    x"3",
        x"5",    x"E",    x"6",    x"2",    x"B",    x"9",    x"0",    x"8",
        x"C",    x"3",    x"5",    x"E",    x"6",    x"2",    x"B",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"9",    x"0",    x"C",    x"5",    x"6",    x"B",    x"0",
        x"C",    x"5",    x"6",    x"B",    x"1",    x"D",    x"4",    x"7",
        x"A",    x"1",    x"D",    x"4",    x"7",    x"A",    x"2",    x"E",
        x"3",    x"8",    x"9",    x"2",    x"E",    x"3",    x"8",    x"9",
        x"3",    x"E",    x"2",    x"9",    x"8",    x"3",    x"E",    x"2",
        x"9",    x"8",    x"4",    x"D",    x"1",    x"A",    x"7",    x"4",
        x"D",    x"1",    x"A",    x"7",    x"4",    x"C",    x"0",    x"B",
        x"6",    x"1",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"5",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"4",    x"6",    x"8",    x"9",
        x"B",    x"D",    x"E",    x"D",    x"B",    x"9",    x"7",    x"6",
        x"4",    x"2",    x"0",    x"1",    x"2",    x"4",    x"6",    x"8",
        x"A",    x"B",    x"D",    x"E",    x"C",    x"B",    x"9",    x"7",
        x"5",    x"3",    x"2",    x"0",    x"1",    x"3",    x"4",    x"6",
        x"8",    x"A",    x"C",    x"D",    x"E",    x"C",    x"A",    x"9",
        x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",    x"5",
        x"7",    x"8",    x"A",    x"C",    x"E",    x"E",    x"C",    x"A",
        x"8",    x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",
        x"5",    x"7",    x"9",    x"A",    x"C",    x"E",    x"D",    x"C",
        x"A",    x"8",    x"6",    x"5",    x"6",    x"8",    x"C",    x"C",
        x"8",    x"4",    x"0",    x"4",    x"9",    x"D",    x"B",    x"7",
        x"2",    x"1",    x"6",    x"A",    x"E",    x"A",    x"6",    x"1",
        x"2",    x"7",    x"B",    x"D",    x"9",    x"5",    x"0",    x"3",
        x"8",    x"C",    x"C",    x"8",    x"3",    x"0",    x"5",    x"9",
        x"D",    x"B",    x"7",    x"2",    x"1",    x"6",    x"A",    x"E",
        x"A",    x"6",    x"1",    x"2",    x"7",    x"B",    x"D",    x"9",
        x"4",    x"0",    x"4",    x"8",    x"D",    x"C",    x"8",    x"3",
        x"0",    x"5",    x"9",    x"E",    x"B",    x"6",    x"0",    x"5",
        x"B",    x"C",    x"6",    x"0",    x"5",    x"B",    x"C",    x"6",
        x"0",    x"5",    x"B",    x"C",    x"6",    x"0",    x"6",    x"C",
        x"B",    x"5",    x"0",    x"6",    x"C",    x"B",    x"5",    x"0",
        x"6",    x"C",    x"B",    x"5",    x"0",    x"6",    x"C",    x"B",
        x"5",    x"0",    x"6",    x"C",    x"B",    x"5",    x"0",    x"6",
        x"C",    x"B",    x"5",    x"0",    x"6",    x"C",    x"B",    x"5",
        x"1",    x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",
        x"A",    x"4",    x"1",    x"7",    x"D",    x"A",    x"4",    x"1",
        x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",    x"A",
        x"4",    x"2",    x"C",    x"8",    x"0",    x"9",    x"B",    x"2",
        x"6",    x"E",    x"5",    x"3",    x"C",    x"8",    x"0",    x"9",
        x"B",    x"2",    x"6",    x"F",    x"6",    x"3",    x"C",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"2",    x"B",    x"9",    x"0",    x"8",    x"C",    x"3",
        x"5",    x"E",    x"6",    x"2",    x"B",    x"9",    x"0",    x"8",
        x"C",    x"3",    x"5",    x"E",    x"6",    x"2",    x"B",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"9",    x"0",    x"C",    x"5",    x"6",    x"B",    x"0",
        x"C",    x"5",    x"6",    x"B",    x"1",    x"D",    x"4",    x"7",
        x"A",    x"1",    x"D",    x"4",    x"7",    x"A",    x"2",    x"E",
        x"3",    x"8",    x"9",    x"2",    x"E",    x"3",    x"8",    x"9",
        x"3",    x"E",    x"2",    x"9",    x"8",    x"3",    x"E",    x"2",
        x"9",    x"8",    x"4",    x"D",    x"1",    x"A",    x"7",    x"4",
        x"D",    x"1",    x"A",    x"7",    x"4",    x"C",    x"0",    x"B",
        x"6",    x"1",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"3",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"4",    x"6",    x"8",    x"9",
        x"B",    x"D",    x"E",    x"D",    x"B",    x"9",    x"7",    x"6",
        x"4",    x"2",    x"0",    x"1",    x"2",    x"4",    x"6",    x"8",
        x"A",    x"B",    x"D",    x"E",    x"C",    x"B",    x"9",    x"7",
        x"5",    x"3",    x"2",    x"0",    x"1",    x"3",    x"4",    x"6",
        x"8",    x"A",    x"C",    x"D",    x"E",    x"C",    x"A",    x"9",
        x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",    x"5",
        x"7",    x"8",    x"A",    x"C",    x"E",    x"E",    x"C",    x"A",
        x"8",    x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",
        x"5",    x"7",    x"9",    x"A",    x"C",    x"E",    x"D",    x"C",
        x"A",    x"8",    x"6",    x"5",    x"6",    x"8",    x"C",    x"C",
        x"8",    x"4",    x"0",    x"4",    x"9",    x"D",    x"B",    x"7",
        x"2",    x"1",    x"6",    x"A",    x"E",    x"A",    x"6",    x"1",
        x"2",    x"7",    x"B",    x"D",    x"9",    x"5",    x"0",    x"3",
        x"8",    x"C",    x"C",    x"8",    x"3",    x"0",    x"5",    x"9",
        x"D",    x"B",    x"7",    x"2",    x"1",    x"6",    x"A",    x"E",
        x"A",    x"6",    x"1",    x"2",    x"7",    x"B",    x"D",    x"9",
        x"4",    x"0",    x"4",    x"8",    x"D",    x"C",    x"8",    x"3",
        x"0",    x"5",    x"9",    x"E",    x"B",    x"6",    x"0",    x"5",
        x"B",    x"C",    x"6",    x"0",    x"5",    x"B",    x"C",    x"6",
        x"0",    x"5",    x"B",    x"C",    x"6",    x"0",    x"6",    x"C",
        x"B",    x"5",    x"0",    x"6",    x"C",    x"B",    x"5",    x"0",
        x"6",    x"C",    x"B",    x"5",    x"0",    x"6",    x"C",    x"B",
        x"5",    x"0",    x"6",    x"C",    x"B",    x"5",    x"0",    x"6",
        x"C",    x"B",    x"5",    x"0",    x"6",    x"C",    x"B",    x"5",
        x"1",    x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",
        x"A",    x"4",    x"1",    x"7",    x"D",    x"A",    x"4",    x"1",
        x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",    x"A",
        x"4",    x"2",    x"C",    x"8",    x"0",    x"9",    x"B",    x"2",
        x"6",    x"E",    x"5",    x"3",    x"C",    x"8",    x"0",    x"9",
        x"B",    x"2",    x"6",    x"F",    x"6",    x"3",    x"C",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"2",    x"B",    x"9",    x"0",    x"8",    x"C",    x"3",
        x"5",    x"E",    x"6",    x"2",    x"B",    x"9",    x"0",    x"8",
        x"C",    x"3",    x"5",    x"E",    x"6",    x"2",    x"B",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"9",    x"0",    x"C",    x"5",    x"6",    x"B",    x"0",
        x"C",    x"5",    x"6",    x"B",    x"1",    x"D",    x"4",    x"7",
        x"A",    x"1",    x"D",    x"4",    x"7",    x"A",    x"2",    x"E",
        x"3",    x"8",    x"9",    x"2",    x"E",    x"3",    x"8",    x"9",
        x"3",    x"E",    x"2",    x"9",    x"8",    x"3",    x"E",    x"2",
        x"9",    x"8",    x"4",    x"D",    x"1",    x"A",    x"7",    x"4",
        x"D",    x"1",    x"A",    x"7",    x"4",    x"C",    x"0",    x"B",
        x"6",    x"1",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"3",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"6",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"4",    x"6",    x"8",    x"9",
        x"B",    x"D",    x"E",    x"D",    x"B",    x"9",    x"7",    x"6",
        x"4",    x"2",    x"0",    x"1",    x"2",    x"4",    x"6",    x"8",
        x"A",    x"B",    x"D",    x"E",    x"C",    x"B",    x"9",    x"7",
        x"5",    x"3",    x"2",    x"0",    x"1",    x"3",    x"4",    x"6",
        x"8",    x"A",    x"C",    x"D",    x"E",    x"C",    x"A",    x"9",
        x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",    x"5",
        x"7",    x"8",    x"A",    x"C",    x"E",    x"E",    x"C",    x"A",
        x"8",    x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",
        x"5",    x"7",    x"9",    x"A",    x"C",    x"E",    x"D",    x"C",
        x"A",    x"8",    x"6",    x"5",    x"6",    x"8",    x"C",    x"C",
        x"8",    x"4",    x"0",    x"4",    x"9",    x"D",    x"B",    x"7",
        x"2",    x"1",    x"6",    x"A",    x"E",    x"A",    x"6",    x"1",
        x"2",    x"7",    x"B",    x"D",    x"9",    x"5",    x"0",    x"3",
        x"8",    x"C",    x"C",    x"8",    x"3",    x"0",    x"5",    x"9",
        x"D",    x"B",    x"7",    x"2",    x"1",    x"6",    x"A",    x"E",
        x"A",    x"6",    x"1",    x"2",    x"7",    x"B",    x"D",    x"9",
        x"4",    x"0",    x"4",    x"8",    x"D",    x"C",    x"8",    x"3",
        x"0",    x"5",    x"9",    x"E",    x"B",    x"6",    x"0",    x"5",
        x"B",    x"C",    x"6",    x"0",    x"5",    x"B",    x"C",    x"6",
        x"0",    x"5",    x"B",    x"C",    x"6",    x"0",    x"6",    x"C",
        x"B",    x"5",    x"0",    x"6",    x"C",    x"B",    x"5",    x"0",
        x"6",    x"C",    x"B",    x"5",    x"0",    x"6",    x"C",    x"B",
        x"5",    x"0",    x"6",    x"C",    x"B",    x"5",    x"0",    x"6",
        x"C",    x"B",    x"5",    x"0",    x"6",    x"C",    x"B",    x"5",
        x"1",    x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",
        x"A",    x"4",    x"1",    x"7",    x"D",    x"A",    x"4",    x"1",
        x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",    x"A",
        x"4",    x"2",    x"C",    x"8",    x"0",    x"9",    x"B",    x"2",
        x"6",    x"E",    x"5",    x"3",    x"C",    x"8",    x"0",    x"9",
        x"B",    x"2",    x"6",    x"F",    x"6",    x"3",    x"C",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"2",    x"B",    x"9",    x"0",    x"8",    x"C",    x"3",
        x"5",    x"E",    x"6",    x"2",    x"B",    x"9",    x"0",    x"8",
        x"C",    x"3",    x"5",    x"E",    x"6",    x"2",    x"B",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"9",    x"0",    x"C",    x"5",    x"6",    x"B",    x"0",
        x"C",    x"5",    x"6",    x"B",    x"1",    x"D",    x"4",    x"7",
        x"A",    x"1",    x"D",    x"4",    x"7",    x"A",    x"2",    x"E",
        x"3",    x"8",    x"9",    x"2",    x"E",    x"3",    x"8",    x"9",
        x"3",    x"E",    x"2",    x"9",    x"8",    x"3",    x"E",    x"2",
        x"9",    x"8",    x"4",    x"D",    x"1",    x"A",    x"7",    x"4",
        x"D",    x"1",    x"A",    x"7",    x"4",    x"C",    x"0",    x"B",
        x"6",    x"1",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"6",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"4",    x"6",    x"8",    x"9",
        x"B",    x"D",    x"E",    x"D",    x"B",    x"9",    x"7",    x"6",
        x"4",    x"2",    x"0",    x"1",    x"2",    x"4",    x"6",    x"8",
        x"A",    x"B",    x"D",    x"E",    x"C",    x"B",    x"9",    x"7",
        x"5",    x"3",    x"2",    x"0",    x"1",    x"3",    x"4",    x"6",
        x"8",    x"A",    x"C",    x"D",    x"E",    x"C",    x"A",    x"9",
        x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",    x"5",
        x"7",    x"8",    x"A",    x"C",    x"E",    x"E",    x"C",    x"A",
        x"8",    x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",
        x"5",    x"7",    x"9",    x"A",    x"C",    x"E",    x"D",    x"C",
        x"A",    x"8",    x"6",    x"5",    x"6",    x"8",    x"C",    x"C",
        x"8",    x"4",    x"0",    x"4",    x"9",    x"D",    x"B",    x"7",
        x"2",    x"1",    x"6",    x"A",    x"E",    x"A",    x"6",    x"1",
        x"2",    x"7",    x"B",    x"D",    x"9",    x"5",    x"0",    x"3",
        x"8",    x"C",    x"C",    x"8",    x"3",    x"0",    x"5",    x"9",
        x"D",    x"B",    x"7",    x"2",    x"1",    x"6",    x"A",    x"E",
        x"A",    x"6",    x"1",    x"2",    x"7",    x"B",    x"D",    x"9",
        x"4",    x"0",    x"4",    x"8",    x"D",    x"C",    x"8",    x"3",
        x"0",    x"5",    x"9",    x"E",    x"B",    x"6",    x"0",    x"5",
        x"B",    x"C",    x"6",    x"0",    x"5",    x"B",    x"C",    x"6",
        x"0",    x"5",    x"B",    x"C",    x"6",    x"0",    x"6",    x"C",
        x"B",    x"5",    x"0",    x"6",    x"C",    x"B",    x"5",    x"0",
        x"6",    x"C",    x"B",    x"5",    x"0",    x"6",    x"C",    x"B",
        x"5",    x"0",    x"6",    x"C",    x"B",    x"5",    x"0",    x"6",
        x"C",    x"B",    x"5",    x"0",    x"6",    x"C",    x"B",    x"5",
        x"1",    x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",
        x"A",    x"4",    x"1",    x"7",    x"D",    x"A",    x"4",    x"1",
        x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",    x"A",
        x"4",    x"2",    x"C",    x"8",    x"0",    x"9",    x"B",    x"2",
        x"6",    x"E",    x"5",    x"3",    x"C",    x"8",    x"0",    x"9",
        x"B",    x"2",    x"6",    x"F",    x"6",    x"3",    x"C",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"2",    x"B",    x"9",    x"0",    x"8",    x"C",    x"3",
        x"5",    x"E",    x"6",    x"2",    x"B",    x"9",    x"0",    x"8",
        x"C",    x"3",    x"5",    x"E",    x"6",    x"2",    x"B",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"9",    x"0",    x"C",    x"5",    x"6",    x"B",    x"0",
        x"C",    x"5",    x"6",    x"B",    x"1",    x"D",    x"4",    x"7",
        x"A",    x"1",    x"D",    x"4",    x"7",    x"A",    x"2",    x"E",
        x"3",    x"8",    x"9",    x"2",    x"E",    x"3",    x"8",    x"9",
        x"3",    x"E",    x"2",    x"9",    x"8",    x"3",    x"E",    x"2",
        x"9",    x"8",    x"4",    x"D",    x"1",    x"A",    x"7",    x"4",
        x"D",    x"1",    x"A",    x"7",    x"4",    x"C",    x"0",    x"B",
        x"6",    x"1",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"5",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"4",    x"6",    x"8",    x"9",
        x"B",    x"D",    x"E",    x"D",    x"B",    x"9",    x"7",    x"6",
        x"4",    x"2",    x"0",    x"1",    x"2",    x"4",    x"6",    x"8",
        x"A",    x"B",    x"D",    x"E",    x"C",    x"B",    x"9",    x"7",
        x"5",    x"3",    x"2",    x"0",    x"1",    x"3",    x"4",    x"6",
        x"8",    x"A",    x"C",    x"D",    x"E",    x"C",    x"A",    x"9",
        x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",    x"5",
        x"7",    x"8",    x"A",    x"C",    x"E",    x"E",    x"C",    x"A",
        x"8",    x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",
        x"5",    x"7",    x"9",    x"A",    x"C",    x"E",    x"D",    x"C",
        x"A",    x"8",    x"6",    x"5",    x"6",    x"8",    x"C",    x"C",
        x"8",    x"4",    x"0",    x"4",    x"9",    x"D",    x"B",    x"7",
        x"2",    x"1",    x"6",    x"A",    x"E",    x"A",    x"6",    x"1",
        x"2",    x"7",    x"B",    x"D",    x"9",    x"5",    x"0",    x"3",
        x"8",    x"C",    x"C",    x"8",    x"3",    x"0",    x"5",    x"9",
        x"D",    x"B",    x"7",    x"2",    x"1",    x"6",    x"A",    x"E",
        x"A",    x"6",    x"1",    x"2",    x"7",    x"B",    x"D",    x"9",
        x"4",    x"0",    x"4",    x"8",    x"D",    x"C",    x"8",    x"3",
        x"0",    x"5",    x"9",    x"E",    x"B",    x"6",    x"0",    x"5",
        x"B",    x"C",    x"6",    x"0",    x"5",    x"B",    x"C",    x"6",
        x"0",    x"5",    x"B",    x"C",    x"6",    x"0",    x"6",    x"C",
        x"B",    x"5",    x"0",    x"6",    x"C",    x"B",    x"5",    x"0",
        x"6",    x"C",    x"B",    x"5",    x"0",    x"6",    x"C",    x"B",
        x"5",    x"0",    x"6",    x"C",    x"B",    x"5",    x"0",    x"6",
        x"C",    x"B",    x"5",    x"0",    x"6",    x"C",    x"B",    x"5",
        x"1",    x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",
        x"A",    x"4",    x"1",    x"7",    x"D",    x"A",    x"4",    x"1",
        x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",    x"A",
        x"4",    x"2",    x"C",    x"8",    x"0",    x"9",    x"B",    x"2",
        x"6",    x"E",    x"5",    x"3",    x"C",    x"8",    x"0",    x"9",
        x"B",    x"2",    x"6",    x"F",    x"6",    x"3",    x"C",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"2",    x"B",    x"9",    x"0",    x"8",    x"C",    x"3",
        x"5",    x"E",    x"6",    x"2",    x"B",    x"9",    x"0",    x"8",
        x"C",    x"3",    x"5",    x"E",    x"6",    x"2",    x"B",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"9",    x"0",    x"C",    x"5",    x"6",    x"B",    x"0",
        x"C",    x"5",    x"6",    x"B",    x"1",    x"D",    x"4",    x"7",
        x"A",    x"1",    x"D",    x"4",    x"7",    x"A",    x"2",    x"E",
        x"3",    x"8",    x"9",    x"2",    x"E",    x"3",    x"8",    x"9",
        x"3",    x"E",    x"2",    x"9",    x"8",    x"3",    x"E",    x"2",
        x"9",    x"8",    x"4",    x"D",    x"1",    x"A",    x"7",    x"4",
        x"D",    x"1",    x"A",    x"7",    x"4",    x"C",    x"0",    x"B",
        x"6",    x"1",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"5",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"4",    x"6",    x"8",    x"9",
        x"B",    x"D",    x"E",    x"D",    x"B",    x"9",    x"7",    x"6",
        x"4",    x"2",    x"0",    x"1",    x"2",    x"4",    x"6",    x"8",
        x"A",    x"B",    x"D",    x"E",    x"C",    x"B",    x"9",    x"7",
        x"5",    x"3",    x"2",    x"0",    x"1",    x"3",    x"4",    x"6",
        x"8",    x"A",    x"C",    x"D",    x"E",    x"C",    x"A",    x"9",
        x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",    x"5",
        x"7",    x"8",    x"A",    x"C",    x"E",    x"E",    x"C",    x"A",
        x"8",    x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",
        x"5",    x"7",    x"9",    x"A",    x"C",    x"E",    x"D",    x"C",
        x"A",    x"8",    x"6",    x"5",    x"6",    x"8",    x"C",    x"C",
        x"8",    x"4",    x"0",    x"4",    x"9",    x"D",    x"B",    x"7",
        x"2",    x"1",    x"6",    x"A",    x"E",    x"A",    x"6",    x"1",
        x"2",    x"7",    x"B",    x"D",    x"9",    x"5",    x"0",    x"3",
        x"8",    x"C",    x"C",    x"8",    x"3",    x"0",    x"5",    x"9",
        x"D",    x"B",    x"7",    x"2",    x"1",    x"6",    x"A",    x"E",
        x"A",    x"6",    x"1",    x"2",    x"7",    x"B",    x"D",    x"9",
        x"4",    x"0",    x"4",    x"8",    x"D",    x"C",    x"8",    x"3",
        x"0",    x"5",    x"9",    x"E",    x"B",    x"6",    x"0",    x"5",
        x"B",    x"C",    x"6",    x"0",    x"5",    x"B",    x"C",    x"6",
        x"0",    x"5",    x"B",    x"C",    x"6",    x"0",    x"6",    x"C",
        x"B",    x"5",    x"0",    x"6",    x"C",    x"B",    x"5",    x"0",
        x"6",    x"C",    x"B",    x"5",    x"0",    x"6",    x"C",    x"B",
        x"5",    x"0",    x"6",    x"C",    x"B",    x"5",    x"0",    x"6",
        x"C",    x"B",    x"5",    x"0",    x"6",    x"C",    x"B",    x"5",
        x"1",    x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",
        x"A",    x"4",    x"1",    x"7",    x"D",    x"A",    x"4",    x"1",
        x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",    x"A",
        x"4",    x"2",    x"C",    x"8",    x"0",    x"9",    x"B",    x"2",
        x"6",    x"E",    x"5",    x"3",    x"C",    x"8",    x"0",    x"9",
        x"B",    x"2",    x"6",    x"F",    x"6",    x"3",    x"C",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"2",    x"B",    x"9",    x"0",    x"8",    x"C",    x"3",
        x"5",    x"E",    x"6",    x"2",    x"B",    x"9",    x"0",    x"8",
        x"C",    x"3",    x"5",    x"E",    x"6",    x"2",    x"B",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"9",    x"0",    x"C",    x"5",    x"6",    x"B",    x"0",
        x"C",    x"5",    x"6",    x"B",    x"1",    x"D",    x"4",    x"7",
        x"A",    x"1",    x"D",    x"4",    x"7",    x"A",    x"2",    x"E",
        x"3",    x"8",    x"9",    x"2",    x"E",    x"3",    x"8",    x"9",
        x"3",    x"E",    x"2",    x"9",    x"8",    x"3",    x"E",    x"2",
        x"9",    x"8",    x"4",    x"D",    x"1",    x"A",    x"7",    x"4",
        x"D",    x"1",    x"A",    x"7",    x"4",    x"C",    x"0",    x"B",
        x"6",    x"1",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"4",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"4",    x"6",    x"8",    x"9",
        x"B",    x"D",    x"E",    x"D",    x"B",    x"9",    x"7",    x"6",
        x"4",    x"2",    x"0",    x"1",    x"2",    x"4",    x"6",    x"8",
        x"A",    x"B",    x"D",    x"E",    x"C",    x"B",    x"9",    x"7",
        x"5",    x"3",    x"2",    x"0",    x"1",    x"3",    x"4",    x"6",
        x"8",    x"A",    x"C",    x"D",    x"E",    x"C",    x"A",    x"9",
        x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",    x"5",
        x"7",    x"8",    x"A",    x"C",    x"E",    x"E",    x"C",    x"A",
        x"8",    x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",
        x"5",    x"7",    x"9",    x"A",    x"C",    x"E",    x"D",    x"C",
        x"A",    x"8",    x"6",    x"5",    x"6",    x"8",    x"C",    x"C",
        x"8",    x"4",    x"0",    x"4",    x"9",    x"D",    x"B",    x"7",
        x"2",    x"1",    x"6",    x"A",    x"E",    x"A",    x"6",    x"1",
        x"2",    x"7",    x"B",    x"D",    x"9",    x"5",    x"0",    x"3",
        x"8",    x"C",    x"C",    x"8",    x"3",    x"0",    x"5",    x"9",
        x"D",    x"B",    x"7",    x"2",    x"1",    x"6",    x"A",    x"E",
        x"A",    x"6",    x"1",    x"2",    x"7",    x"B",    x"D",    x"9",
        x"4",    x"0",    x"4",    x"8",    x"D",    x"C",    x"8",    x"3",
        x"0",    x"5",    x"9",    x"E",    x"B",    x"6",    x"0",    x"5",
        x"B",    x"C",    x"6",    x"0",    x"5",    x"B",    x"C",    x"6",
        x"0",    x"5",    x"B",    x"C",    x"6",    x"0",    x"6",    x"C",
        x"B",    x"5",    x"0",    x"6",    x"C",    x"B",    x"5",    x"0",
        x"6",    x"C",    x"B",    x"5",    x"0",    x"6",    x"C",    x"B",
        x"5",    x"0",    x"6",    x"C",    x"B",    x"5",    x"0",    x"6",
        x"C",    x"B",    x"5",    x"0",    x"6",    x"C",    x"B",    x"5",
        x"1",    x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",
        x"A",    x"4",    x"1",    x"7",    x"D",    x"A",    x"4",    x"1",
        x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",    x"A",
        x"4",    x"2",    x"C",    x"8",    x"0",    x"9",    x"B",    x"2",
        x"6",    x"E",    x"5",    x"3",    x"C",    x"8",    x"0",    x"9",
        x"B",    x"2",    x"6",    x"F",    x"6",    x"3",    x"C",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"2",    x"B",    x"9",    x"0",    x"8",    x"C",    x"3",
        x"5",    x"E",    x"6",    x"2",    x"B",    x"9",    x"0",    x"8",
        x"C",    x"3",    x"5",    x"E",    x"6",    x"2",    x"B",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"9",    x"0",    x"C",    x"5",    x"6",    x"B",    x"0",
        x"C",    x"5",    x"6",    x"B",    x"1",    x"D",    x"4",    x"7",
        x"A",    x"1",    x"D",    x"4",    x"7",    x"A",    x"2",    x"E",
        x"3",    x"8",    x"9",    x"2",    x"E",    x"3",    x"8",    x"9",
        x"3",    x"E",    x"2",    x"9",    x"8",    x"3",    x"E",    x"2",
        x"9",    x"8",    x"4",    x"D",    x"1",    x"A",    x"7",    x"4",
        x"D",    x"1",    x"A",    x"7",    x"4",    x"C",    x"0",    x"B",
        x"6",    x"1",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"4",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"8",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"4",    x"6",    x"8",    x"9",
        x"B",    x"D",    x"E",    x"D",    x"B",    x"9",    x"7",    x"6",
        x"4",    x"2",    x"0",    x"1",    x"2",    x"4",    x"6",    x"8",
        x"A",    x"B",    x"D",    x"E",    x"C",    x"B",    x"9",    x"7",
        x"5",    x"3",    x"2",    x"0",    x"1",    x"3",    x"4",    x"6",
        x"8",    x"A",    x"C",    x"D",    x"E",    x"C",    x"A",    x"9",
        x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",    x"5",
        x"7",    x"8",    x"A",    x"C",    x"E",    x"E",    x"C",    x"A",
        x"8",    x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",
        x"5",    x"7",    x"9",    x"A",    x"C",    x"E",    x"D",    x"C",
        x"A",    x"8",    x"6",    x"5",    x"6",    x"8",    x"C",    x"C",
        x"8",    x"4",    x"0",    x"4",    x"9",    x"D",    x"B",    x"7",
        x"2",    x"1",    x"6",    x"A",    x"E",    x"A",    x"6",    x"1",
        x"2",    x"7",    x"B",    x"D",    x"9",    x"5",    x"0",    x"3",
        x"8",    x"C",    x"C",    x"8",    x"3",    x"0",    x"5",    x"9",
        x"D",    x"B",    x"7",    x"2",    x"1",    x"6",    x"A",    x"E",
        x"A",    x"6",    x"1",    x"2",    x"7",    x"B",    x"D",    x"9",
        x"4",    x"0",    x"4",    x"8",    x"D",    x"C",    x"8",    x"3",
        x"0",    x"5",    x"9",    x"E",    x"B",    x"6",    x"0",    x"5",
        x"B",    x"C",    x"6",    x"0",    x"5",    x"B",    x"C",    x"6",
        x"0",    x"5",    x"B",    x"C",    x"6",    x"0",    x"6",    x"C",
        x"B",    x"5",    x"0",    x"6",    x"C",    x"B",    x"5",    x"0",
        x"6",    x"C",    x"B",    x"5",    x"0",    x"6",    x"C",    x"B",
        x"5",    x"0",    x"6",    x"C",    x"B",    x"5",    x"0",    x"6",
        x"C",    x"B",    x"5",    x"0",    x"6",    x"C",    x"B",    x"5",
        x"1",    x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",
        x"A",    x"4",    x"1",    x"7",    x"D",    x"A",    x"4",    x"1",
        x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",    x"A",
        x"4",    x"2",    x"C",    x"8",    x"0",    x"9",    x"B",    x"2",
        x"6",    x"E",    x"5",    x"3",    x"C",    x"8",    x"0",    x"9",
        x"B",    x"2",    x"6",    x"F",    x"6",    x"3",    x"C",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"2",    x"B",    x"9",    x"0",    x"8",    x"C",    x"3",
        x"5",    x"E",    x"6",    x"2",    x"B",    x"9",    x"0",    x"8",
        x"C",    x"3",    x"5",    x"E",    x"6",    x"2",    x"B",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"9",    x"0",    x"C",    x"5",    x"6",    x"B",    x"0",
        x"C",    x"5",    x"6",    x"B",    x"1",    x"D",    x"4",    x"7",
        x"A",    x"1",    x"D",    x"4",    x"7",    x"A",    x"2",    x"E",
        x"3",    x"8",    x"9",    x"2",    x"E",    x"3",    x"8",    x"9",
        x"3",    x"E",    x"2",    x"9",    x"8",    x"3",    x"E",    x"2",
        x"9",    x"8",    x"4",    x"D",    x"1",    x"A",    x"7",    x"4",
        x"D",    x"1",    x"A",    x"7",    x"4",    x"C",    x"0",    x"B",
        x"6",    x"1",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"8",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"E",    x"F",
        x"E",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"D",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"D",    x"3",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"4",    x"6",    x"8",    x"9",
        x"B",    x"D",    x"E",    x"D",    x"B",    x"9",    x"7",    x"6",
        x"4",    x"2",    x"0",    x"1",    x"2",    x"4",    x"6",    x"8",
        x"A",    x"B",    x"D",    x"E",    x"C",    x"B",    x"9",    x"7",
        x"5",    x"3",    x"2",    x"0",    x"1",    x"3",    x"4",    x"6",
        x"8",    x"A",    x"C",    x"D",    x"E",    x"C",    x"A",    x"9",
        x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",    x"5",
        x"7",    x"8",    x"A",    x"C",    x"E",    x"E",    x"C",    x"A",
        x"8",    x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",
        x"5",    x"7",    x"9",    x"A",    x"C",    x"E",    x"D",    x"C",
        x"A",    x"8",    x"6",    x"5",    x"6",    x"8",    x"C",    x"C",
        x"8",    x"4",    x"0",    x"4",    x"9",    x"D",    x"B",    x"7",
        x"2",    x"1",    x"6",    x"A",    x"E",    x"A",    x"6",    x"1",
        x"2",    x"7",    x"B",    x"D",    x"9",    x"5",    x"0",    x"3",
        x"8",    x"C",    x"C",    x"8",    x"3",    x"0",    x"5",    x"9",
        x"D",    x"B",    x"7",    x"2",    x"1",    x"6",    x"A",    x"E",
        x"A",    x"6",    x"1",    x"2",    x"7",    x"B",    x"D",    x"9",
        x"4",    x"0",    x"4",    x"8",    x"D",    x"C",    x"8",    x"3",
        x"0",    x"5",    x"9",    x"E",    x"B",    x"6",    x"0",    x"5",
        x"B",    x"C",    x"6",    x"0",    x"5",    x"B",    x"C",    x"6",
        x"0",    x"5",    x"B",    x"C",    x"6",    x"0",    x"6",    x"C",
        x"B",    x"5",    x"0",    x"6",    x"C",    x"B",    x"5",    x"0",
        x"6",    x"C",    x"B",    x"5",    x"0",    x"6",    x"C",    x"B",
        x"5",    x"0",    x"6",    x"C",    x"B",    x"5",    x"0",    x"6",
        x"C",    x"B",    x"5",    x"0",    x"6",    x"C",    x"B",    x"5",
        x"1",    x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",
        x"A",    x"4",    x"1",    x"7",    x"D",    x"A",    x"4",    x"1",
        x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",    x"A",
        x"4",    x"2",    x"C",    x"8",    x"0",    x"9",    x"B",    x"2",
        x"6",    x"E",    x"5",    x"3",    x"C",    x"8",    x"0",    x"9",
        x"B",    x"2",    x"6",    x"F",    x"6",    x"3",    x"C",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"2",    x"B",    x"9",    x"0",    x"8",    x"C",    x"3",
        x"5",    x"E",    x"6",    x"2",    x"B",    x"9",    x"0",    x"8",
        x"C",    x"3",    x"5",    x"E",    x"6",    x"2",    x"B",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"9",    x"0",    x"C",    x"5",    x"6",    x"B",    x"0",
        x"C",    x"5",    x"6",    x"B",    x"1",    x"D",    x"4",    x"7",
        x"A",    x"1",    x"D",    x"4",    x"7",    x"A",    x"2",    x"E",
        x"3",    x"8",    x"9",    x"2",    x"E",    x"3",    x"8",    x"9",
        x"3",    x"E",    x"2",    x"9",    x"8",    x"3",    x"E",    x"2",
        x"9",    x"8",    x"4",    x"D",    x"1",    x"A",    x"7",    x"4",
        x"D",    x"1",    x"A",    x"7",    x"4",    x"C",    x"0",    x"B",
        x"6",    x"1",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"3",    x"D",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"D",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"E",
        x"F",    x"E",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"A",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"2",    x"4",    x"6",    x"8",    x"9",
        x"B",    x"D",    x"E",    x"D",    x"B",    x"9",    x"7",    x"6",
        x"4",    x"2",    x"0",    x"1",    x"2",    x"4",    x"6",    x"8",
        x"A",    x"B",    x"D",    x"E",    x"C",    x"B",    x"9",    x"7",
        x"5",    x"3",    x"2",    x"0",    x"1",    x"3",    x"4",    x"6",
        x"8",    x"A",    x"C",    x"D",    x"E",    x"C",    x"A",    x"9",
        x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",    x"5",
        x"7",    x"8",    x"A",    x"C",    x"E",    x"E",    x"C",    x"A",
        x"8",    x"7",    x"5",    x"3",    x"1",    x"0",    x"1",    x"3",
        x"5",    x"7",    x"9",    x"A",    x"C",    x"E",    x"D",    x"C",
        x"A",    x"8",    x"6",    x"5",    x"6",    x"8",    x"C",    x"C",
        x"8",    x"4",    x"0",    x"4",    x"9",    x"D",    x"B",    x"7",
        x"2",    x"1",    x"6",    x"A",    x"E",    x"A",    x"6",    x"1",
        x"2",    x"7",    x"B",    x"D",    x"9",    x"5",    x"0",    x"3",
        x"8",    x"C",    x"C",    x"8",    x"3",    x"0",    x"5",    x"9",
        x"D",    x"B",    x"7",    x"2",    x"1",    x"6",    x"A",    x"E",
        x"A",    x"6",    x"1",    x"2",    x"7",    x"B",    x"D",    x"9",
        x"4",    x"0",    x"4",    x"8",    x"D",    x"C",    x"8",    x"3",
        x"0",    x"5",    x"9",    x"E",    x"B",    x"6",    x"0",    x"5",
        x"B",    x"C",    x"6",    x"0",    x"5",    x"B",    x"C",    x"6",
        x"0",    x"5",    x"B",    x"C",    x"6",    x"0",    x"6",    x"C",
        x"B",    x"5",    x"0",    x"6",    x"C",    x"B",    x"5",    x"0",
        x"6",    x"C",    x"B",    x"5",    x"0",    x"6",    x"C",    x"B",
        x"5",    x"0",    x"6",    x"C",    x"B",    x"5",    x"0",    x"6",
        x"C",    x"B",    x"5",    x"0",    x"6",    x"C",    x"B",    x"5",
        x"1",    x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",
        x"A",    x"4",    x"1",    x"7",    x"D",    x"A",    x"4",    x"1",
        x"7",    x"D",    x"A",    x"4",    x"1",    x"7",    x"D",    x"A",
        x"4",    x"2",    x"C",    x"8",    x"0",    x"9",    x"B",    x"2",
        x"6",    x"E",    x"5",    x"3",    x"C",    x"8",    x"0",    x"9",
        x"B",    x"2",    x"6",    x"F",    x"6",    x"3",    x"C",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"2",    x"B",    x"9",    x"0",    x"8",    x"C",    x"3",
        x"5",    x"E",    x"6",    x"2",    x"B",    x"9",    x"0",    x"8",
        x"C",    x"3",    x"5",    x"E",    x"6",    x"2",    x"B",    x"9",
        x"0",    x"8",    x"C",    x"3",    x"5",    x"E",    x"6",    x"2",
        x"B",    x"9",    x"0",    x"8",    x"C",    x"3",    x"5",    x"E",
        x"6",    x"9",    x"0",    x"C",    x"5",    x"6",    x"B",    x"0",
        x"C",    x"5",    x"6",    x"B",    x"1",    x"D",    x"4",    x"7",
        x"A",    x"1",    x"D",    x"4",    x"7",    x"A",    x"2",    x"E",
        x"3",    x"8",    x"9",    x"2",    x"E",    x"3",    x"8",    x"9",
        x"3",    x"E",    x"2",    x"9",    x"8",    x"3",    x"E",    x"2",
        x"9",    x"8",    x"4",    x"D",    x"1",    x"A",    x"7",    x"4",
        x"D",    x"1",    x"A",    x"7",    x"4",    x"C",    x"0",    x"B",
        x"6",    x"1",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"A",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"E",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"E",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"E",    x"E",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"2",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"5",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"E",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"D",    x"E",    x"E",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"E",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"E",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"5",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"2",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"5",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"B",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"E",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"B",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"E",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"2",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"5",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"B",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"E",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"E",    x"E",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"5",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"5",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"B",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"E",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"D",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"5",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"B",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"E",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"9",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"5",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"5",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"B",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"E",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"D",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"1",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"5",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"B",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"E",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"E",    x"8",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"5",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"5",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"B",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"E",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"C",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"1",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"5",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"B",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"E",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"E",    x"8",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"5",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"5",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"B",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"E",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"1",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"5",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"B",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"E",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"E",
        x"8",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"6",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"5",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"B",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"E",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"C",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"1",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"5",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"B",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"E",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"E",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"6",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"5",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"B",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"E",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"2",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"5",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"B",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"E",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"E",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"5",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"B",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"E",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"A",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"4",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"5",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"B",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"E",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"E",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"5",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"B",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"E",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"9",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"5",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"5",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"B",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"E",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"1",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"5",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"B",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"E",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"E",    x"8",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"6",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"5",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"B",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"E",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"2",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"5",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"B",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"E",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"E",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"5",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"B",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"E",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"5",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"5",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"B",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"E",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"D",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"1",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"5",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"B",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"E",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"E",
        x"8",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"6",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"5",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"B",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"E",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"B",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"4",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"5",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"B",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"E",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"D",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"1",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"5",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"B",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"E",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"E",    x"8",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"6",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"5",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"B",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"E",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"B",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"5",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"B",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"E",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"E",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"5",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"B",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"E",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"9",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"6",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"5",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"B",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"E",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"C",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"3",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"5",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"B",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"E",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"E",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"1",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"5",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"B",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"E",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"E",    x"8",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"E",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"E",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"E",    x"F",    x"F",    x"E",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"A",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"5",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"B",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"E",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"E",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"E",    x"F",    x"F",    x"E",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"E",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"E",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"7",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"7",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"4",    x"2",    x"2",    x"2",    x"2",    x"2",
        x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",
        x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",
        x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",
        x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",
        x"3",    x"5",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",    x"6",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"9",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"C",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"E",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"A",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"E",    x"F",
        x"E",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"D",    x"F",    x"F",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"E",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"E",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"A",    x"C",    x"C",
        x"6",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"E",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"F",    x"F",    x"D",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"E",
        x"F",    x"E",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"8",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"9",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"E",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"F",
        x"7",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"9",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"8",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"8",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"E",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"F",
        x"7",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"8",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"8",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"E",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"E",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"F",
        x"7",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"E",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"8",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"8",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"8",    x"E",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"E",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"F",
        x"7",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"E",    x"8",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"8",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"8",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"A",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"E",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"F",
        x"7",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"A",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"8",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"8",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"E",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"F",
        x"7",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"C",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"8",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"8",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"E",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"F",
        x"7",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"8",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"8",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"E",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"E",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"F",
        x"7",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"E",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"8",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"8",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"E",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"E",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"F",
        x"7",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"E",    x"9",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"8",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"8",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"E",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"F",
        x"7",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"8",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"8",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"E",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"F",
        x"7",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"8",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"8",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"D",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"E",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"F",
        x"7",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"D",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"8",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"8",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"E",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"E",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"F",
        x"7",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"E",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"8",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"8",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"8",    x"E",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"E",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"F",
        x"7",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"E",    x"8",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"8",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"8",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"9",    x"E",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"E",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"F",
        x"7",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"E",    x"9",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"8",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"8",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"9",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"E",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"F",
        x"7",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"A",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"8",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"8",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"E",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"F",
        x"7",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"8",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"8",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"E",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"F",
        x"7",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"8",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"8",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"E",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"F",
        x"7",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"8",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"8",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"D",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"E",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"F",
        x"7",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"D",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"8",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"8",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"D",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"E",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"F",
        x"7",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"E",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"8",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"8",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"E",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"E",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"F",
        x"7",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"E",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"8",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"8",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"E",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"E",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"F",
        x"7",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"E",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"8",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"8",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"8",    x"E",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"E",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"F",
        x"7",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"E",    x"8",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"8",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"8",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"8",    x"E",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"E",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"F",
        x"7",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"E",    x"8",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"8",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"8",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"E",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"E",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"F",
        x"7",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"E",    x"8",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"8",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"8",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"E",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"E",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"F",
        x"7",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"E",    x"8",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"8",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"8",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"8",
        x"E",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"E",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"F",
        x"7",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"E",
        x"8",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"8",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"8",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"8",    x"E",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"E",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"F",
        x"7",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"E",    x"8",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"8",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"8",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"E",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"E",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"F",
        x"7",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"E",    x"8",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"8",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"8",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"D",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"D",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"F",
        x"7",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"B",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"D",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"8",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"8",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"C",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"D",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"F",
        x"7",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"B",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"C",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"8",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"8",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"C",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"D",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"F",
        x"7",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"B",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"C",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"8",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"8",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"E",    x"D",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"D",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",    x"F",
        x"7",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"B",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"D",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"8",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"8",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"D",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"B",    x"2",    x"2",    x"2",    x"2",    x"2",
        x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",
        x"2",    x"2",    x"2",    x"2",    x"2",    x"C",    x"F",    x"F",
        x"8",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",
        x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",
        x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",
        x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",
        x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",
        x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",
        x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",
        x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",
        x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"1",    x"1",
        x"1",    x"1",    x"1",    x"1",    x"1",    x"1",    x"1",    x"1",
        x"1",    x"1",    x"1",    x"1",    x"1",    x"1",    x"1",    x"1",
        x"1",    x"1",    x"1",    x"1",    x"1",    x"1",    x"1",    x"1",
        x"1",    x"1",    x"1",    x"1",    x"1",    x"1",    x"1",    x"1",
        x"1",    x"1",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",
        x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",
        x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",
        x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",
        x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",
        x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",
        x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",
        x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",
        x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",
        x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",
        x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",
        x"2",    x"2",    x"2",    x"2",    x"2",    x"A",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"D",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"8",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"D",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"8",    x"F",    x"F",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"D",    x"F",    x"F",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"F",    x"F",    x"D",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"F",    x"F",    x"8",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"D",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"8",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"8",    x"8",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"8",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"8",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"8",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"8",    x"8",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"8",    x"8",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"8",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"8",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"9",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"8",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"8",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"9",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"8",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"8",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"9",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"8",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"8",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"8",
        x"8",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"8",
        x"8",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"8",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"8",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"8",    x"8",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"8",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"8",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"8",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"9",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"8",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"8",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"9",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"9",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"8",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"8",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"8",    x"8",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"8",    x"8",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"8",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"8",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"9",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"8",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"8",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"9",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"9",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"8",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"8",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"8",    x"8",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"8",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"8",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"8",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"A",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"8",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"8",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"C",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"C",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"8",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"8",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"D",    x"8",    x"9",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"9",    x"8",    x"D",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"8",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"8",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"D",    x"7",    x"7",    x"9",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"9",    x"7",    x"7",    x"D",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"8",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"8",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"8",
        x"9",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"9",
        x"8",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"8",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"8",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"9",    x"8",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"9",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"8",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"8",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"9",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"9",    x"8",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"8",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"8",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"8",    x"8",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"8",    x"8",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"8",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"8",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"9",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"8",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"8",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"8",
        x"8",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"8",
        x"8",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"8",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"8",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"9",    x"8",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"9",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"8",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"8",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"9",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"9",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"8",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"8",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"8",    x"9",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"9",    x"8",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"8",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"8",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"8",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"8",    x"8",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"8",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"8",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"9",    x"8",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"9",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"8",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"8",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"9",    x"8",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"8",    x"9",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"8",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"8",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"9",    x"8",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"8",    x"9",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"8",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"8",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"8",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"8",    x"9",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"8",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"8",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"9",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"9",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"8",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",    x"5",
        x"5",    x"5",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"C",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"C",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"F",    x"F",    x"C",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"9",    x"F",    x"F",    x"9",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"B",    x"F",    x"F",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"C",    x"F",    x"E",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"9",    x"9",    x"8",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"8",    x"9",    x"9",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"E",    x"F",    x"C",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"F",    x"F",    x"B",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"9",    x"F",    x"F",    x"9",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"C",    x"F",    x"F",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",
        x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"8",    x"C",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"E",    x"C",    x"8",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"8",    x"B",    x"E",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"E",    x"D",    x"9",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"9",    x"C",    x"E",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"D",    x"F",
        x"D",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"F",    x"F",    x"C",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"F",    x"F",
        x"B",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"B",    x"F",    x"F",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"C",    x"F",    x"F",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"D",    x"F",    x"E",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"E",    x"F",    x"D",
        x"A",    x"9",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"A",
        x"D",    x"F",    x"E",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"E",    x"F",    x"D",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"F",    x"F",    x"C",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"F",    x"F",    x"B",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"B",
        x"F",    x"F",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"C",    x"F",    x"F",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"D",
        x"F",    x"D",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",
        x"7",    x"7",    x"8",    x"9",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"9",    x"8",    x"7",    x"7",
        x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"8",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"8",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"8",    x"9",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"8",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"8",
        x"9",    x"8",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"9",
        x"8",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"8",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"9",    x"9",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"8",    x"9",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"8",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"8",    x"9",    x"8",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"8",    x"9",    x"8",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"8",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"8",
        x"9",    x"8",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"9",
        x"8",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"8",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"8",    x"9",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"9",    x"8",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"8",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"9",    x"8",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"8",    x"9",    x"8",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"8",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"8",    x"9",    x"8",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"9",    x"8",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"8",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"9",    x"9",    x"8",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"8",    x"9",    x"9",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"8",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"8",
        x"9",    x"9",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"9",    x"9",
        x"8",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"8",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"F",    x"E",    x"B",    x"9",    x"9",    x"8",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"8",    x"9",    x"9",    x"B",    x"E",    x"F",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"8",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"8",
        x"9",    x"9",    x"8",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"9",    x"9",
        x"8",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"8",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"9",    x"9",    x"9",    x"8",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"8",    x"9",    x"9",    x"9",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"8",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"8",    x"9",    x"9",    x"9",    x"8",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"9",    x"9",    x"8",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"8",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"8",
        x"9",    x"9",    x"9",    x"8",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"8",    x"9",    x"9",    x"9",
        x"8",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"8",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"8",
        x"9",    x"9",    x"9",    x"9",    x"8",    x"8",    x"4",    x"4",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",    x"3",
        x"4",    x"4",    x"8",    x"8",    x"9",    x"9",    x"9",    x"9",
        x"8",    x"8",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"8",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",
        x"7",    x"7",    x"7",    x"8",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"6",    x"6",
        x"6",    x"6",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"8",    x"8",    x"7",    x"7",
        x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"8",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"8",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"8",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"8",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"8",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"8",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"8",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"8",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"8",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"8",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"8",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"8",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"8",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"8",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"C",    x"F",
        x"C",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"8",    x"F",    x"F",
        x"A",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"A",    x"F",    x"F",    x"8",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"F",    x"D",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"D",    x"F",    x"C",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"F",    x"F",    x"B",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"8",    x"F",    x"F",    x"A",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"A",
        x"F",    x"F",    x"8",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"B",    x"F",    x"F",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"C",
        x"F",    x"C",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"D",    x"F",
        x"D",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"F",    x"F",    x"C",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"F",    x"F",
        x"B",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"B",    x"F",    x"F",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"C",    x"F",    x"F",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"D",    x"F",    x"E",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"E",    x"F",    x"D",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"F",    x"F",    x"C",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"F",    x"F",    x"B",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"B",    x"F",    x"F",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"C",    x"F",    x"F",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"D",    x"F",    x"E",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"E",    x"F",    x"D",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"F",    x"F",    x"C",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"F",    x"F",    x"B",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"B",
        x"F",    x"F",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"C",    x"F",    x"F",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"D",
        x"F",    x"D",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"A",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",
        x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",
        x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",
        x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",
        x"2",    x"2",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"6",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",
        x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",
        x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",
        x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",
        x"2",    x"6",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",
        x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",
        x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",
        x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",
        x"2",    x"A",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"A",
        x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",
        x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",
        x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",
        x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",
        x"2",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"6",
        x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",
        x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",
        x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",
        x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",
        x"6",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"2",
        x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",
        x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",
        x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",
        x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",
        x"A",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"A",    x"2",
        x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",
        x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",
        x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",
        x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"6",    x"2",
        x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",
        x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",
        x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",
        x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"6",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"2",    x"2",
        x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",
        x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",
        x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",
        x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"2",    x"A",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"A",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"4",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"4",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"A",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"A",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"4",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"A",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"A",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"4",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"A",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"A",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"4",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"4",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"A",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"A",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"4",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"A",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"A",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"4",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"A",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"A",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"4",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"4",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"A",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"A",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"4",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"A",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"A",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"4",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"A",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"A",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"4",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"4",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"A",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"A",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"4",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"A",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"A",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"4",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"A",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"A",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"4",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"4",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"A",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"A",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"4",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"A",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"A",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"4",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"A",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F"
    );

end package ram_init_phillips_pm5544_grayscale;

