----------------------------------------------------------------------------------
-- Company:
-- Engineer:
--
-- Design Name:
-- Module Name: ram_init_smpte_color_bars_tty16 - Behavioral
-- Project Name:
-- Target Devices:
-- Tool Versions: 2021.2
-- Description:
--
-- Dependencies:
--
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
----------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;


package ram_init_smpte_color_bars_tty16 is

    constant FB_WIDTH : integer := 640;
    constant FB_HEIGHT : integer := 480;
    constant FB_PIXELS : integer := FB_WIDTH * FB_HEIGHT;

    constant DATA_WIDTH : integer := 4;
    constant DEPTH : integer := FB_PIXELS;

    subtype addr_t is integer range 0 to DEPTH - 1;
    subtype ram_word_t is std_logic_vector(DATA_WIDTH-1 downto 0);

    type ram_type is array (addr_t) of ram_word_t;

    -- Synthesizable constant RAM content
    constant INIT_RAM : ram_type := (
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"3",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"B",
        x"B",    x"B",    x"B",    x"B",    x"B",    x"B",    x"3",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"2",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",    x"A",
        x"A",    x"A",    x"A",    x"A",    x"A",    x"2",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"1",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",    x"9",
        x"9",    x"9",    x"9",    x"9",    x"5",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"4",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"5",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"4",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"5",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"4",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"5",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"4",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"5",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"4",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"5",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"4",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"5",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"4",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"5",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"4",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"5",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"4",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"5",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"4",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"5",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"4",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"5",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"4",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"5",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"4",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"5",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"4",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"5",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"4",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"5",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"4",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"5",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"4",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"5",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"4",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"5",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"4",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"5",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"4",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"5",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"4",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"5",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"4",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"5",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"4",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"5",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"4",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"5",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"4",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"5",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"4",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"5",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"4",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"5",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"4",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"5",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"4",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"5",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"4",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"5",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"4",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"5",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"4",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"5",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"4",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"5",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"4",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"5",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"4",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"5",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"4",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"5",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"4",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"5",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"4",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"5",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"4",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"5",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",    x"C",
        x"C",    x"C",    x"C",    x"4",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",    x"D",
        x"D",    x"D",    x"5",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"6",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",    x"E",
        x"E",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"8",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",    x"7",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"7",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",    x"F",
        x"F",    x"F",    x"F",    x"F",    x"8",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",
        x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"4",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",
        x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0",    x"0"
    );

end package ram_init_smpte_color_bars_tty16;

